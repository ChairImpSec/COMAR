//
// -----------------------------------------------------------------
// COMPANY : Ruhr University Bochum
// AUTHOR  : AUTHOR  : David Knichel david.knichel@rub.de and Amir Moradi amir.moradi@rub.de 
// DOCUMENT: [Composable Gadgets with Reused Fresh Masks] https://doi.org/10.46586/tches.v2022.i3.114-140
// -----------------------------------------------------------------
//
// Copyright (c) 2022, David Knichel and  Amir Moradi
//
// All rights reserved.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
// ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
// WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
// DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
// DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
// (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
// LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
// ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
// (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
// SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.
//
// Please see LICENSE and README for license and further instructions.
//

module CRAFT ( clk, rst, plaintext, key, ciphertext, done );
  (* AGEMA = "secure" *) input [63:0]  plaintext;
  (* AGEMA = "secure" *) input [127:0] key;
  (* AGEMA = "clock" *)  input clk;
  (* AGEMA = "reset" *)  input rst;

  output [63:0] ciphertext;
  output done;
 
  wire   RoundConstant_4_, RoundConstant_0, done_internal,
         MCInst_XOR_r0_Inst_0_n2, MCInst_XOR_r0_Inst_0_n1,
         MCInst_XOR_r1_Inst_0_n1, MCInst_XOR_r0_Inst_1_n2,
         MCInst_XOR_r0_Inst_1_n1, MCInst_XOR_r1_Inst_1_n1,
         MCInst_XOR_r0_Inst_2_n2, MCInst_XOR_r0_Inst_2_n1,
         MCInst_XOR_r1_Inst_2_n1, MCInst_XOR_r0_Inst_3_n2,
         MCInst_XOR_r0_Inst_3_n1, MCInst_XOR_r1_Inst_3_n1,
         MCInst_XOR_r0_Inst_4_n2, MCInst_XOR_r0_Inst_4_n1,
         MCInst_XOR_r1_Inst_4_n1, MCInst_XOR_r0_Inst_5_n2,
         MCInst_XOR_r0_Inst_5_n1, MCInst_XOR_r1_Inst_5_n1,
         MCInst_XOR_r0_Inst_6_n2, MCInst_XOR_r0_Inst_6_n1,
         MCInst_XOR_r1_Inst_6_n1, MCInst_XOR_r0_Inst_7_n2,
         MCInst_XOR_r0_Inst_7_n1, MCInst_XOR_r1_Inst_7_n1,
         MCInst_XOR_r0_Inst_8_n2, MCInst_XOR_r0_Inst_8_n1,
         MCInst_XOR_r1_Inst_8_n1, MCInst_XOR_r0_Inst_9_n2,
         MCInst_XOR_r0_Inst_9_n1, MCInst_XOR_r1_Inst_9_n1,
         MCInst_XOR_r0_Inst_10_n2, MCInst_XOR_r0_Inst_10_n1,
         MCInst_XOR_r1_Inst_10_n1, MCInst_XOR_r0_Inst_11_n2,
         MCInst_XOR_r0_Inst_11_n1, MCInst_XOR_r1_Inst_11_n1,
         MCInst_XOR_r0_Inst_12_n2, MCInst_XOR_r0_Inst_12_n1,
         MCInst_XOR_r1_Inst_12_n1, MCInst_XOR_r0_Inst_13_n2,
         MCInst_XOR_r0_Inst_13_n1, MCInst_XOR_r1_Inst_13_n1,
         MCInst_XOR_r0_Inst_14_n2, MCInst_XOR_r0_Inst_14_n1,
         MCInst_XOR_r1_Inst_14_n1, MCInst_XOR_r0_Inst_15_n2,
         MCInst_XOR_r0_Inst_15_n1, MCInst_XOR_r1_Inst_15_n1,
         AddKeyXOR1_XORInst_0_0_n1, AddKeyXOR1_XORInst_0_1_n1,
         AddKeyXOR1_XORInst_0_2_n1, AddKeyXOR1_XORInst_0_3_n1,
         AddKeyXOR1_XORInst_1_0_n1, AddKeyXOR1_XORInst_1_1_n1,
         AddKeyXOR1_XORInst_1_2_n1, AddKeyXOR1_XORInst_1_3_n1,
         AddKeyXOR1_XORInst_2_0_n1, AddKeyXOR1_XORInst_2_1_n1,
         AddKeyXOR1_XORInst_2_2_n1, AddKeyXOR1_XORInst_2_3_n1,
         AddKeyXOR1_XORInst_3_0_n1, AddKeyXOR1_XORInst_3_1_n1,
         AddKeyXOR1_XORInst_3_2_n1, AddKeyXOR1_XORInst_3_3_n1,
         AddKeyConstXOR_XORInst_0_0_n2, AddKeyConstXOR_XORInst_0_0_n1,
         AddKeyConstXOR_XORInst_0_1_n2, AddKeyConstXOR_XORInst_0_1_n1,
         AddKeyConstXOR_XORInst_0_2_n2, AddKeyConstXOR_XORInst_0_2_n1,
         AddKeyConstXOR_XORInst_0_3_n2, AddKeyConstXOR_XORInst_0_3_n1,
         AddKeyConstXOR_XORInst_1_0_n2, AddKeyConstXOR_XORInst_1_0_n1,
         AddKeyConstXOR_XORInst_1_1_n2, AddKeyConstXOR_XORInst_1_1_n1,
         AddKeyConstXOR_XORInst_1_2_n2, AddKeyConstXOR_XORInst_1_2_n1,
         AddKeyConstXOR_XORInst_1_3_n2, AddKeyConstXOR_XORInst_1_3_n1,
         AddKeyXOR2_XORInst_0_0_n1, AddKeyXOR2_XORInst_0_1_n1,
         AddKeyXOR2_XORInst_0_2_n1, AddKeyXOR2_XORInst_0_3_n1,
         AddKeyXOR2_XORInst_1_0_n1, AddKeyXOR2_XORInst_1_1_n1,
         AddKeyXOR2_XORInst_1_2_n1, AddKeyXOR2_XORInst_1_3_n1,
         AddKeyXOR2_XORInst_2_0_n1, AddKeyXOR2_XORInst_2_1_n1,
         AddKeyXOR2_XORInst_2_2_n1, AddKeyXOR2_XORInst_2_3_n1,
         AddKeyXOR2_XORInst_3_0_n1, AddKeyXOR2_XORInst_3_1_n1,
         AddKeyXOR2_XORInst_3_2_n1, AddKeyXOR2_XORInst_3_3_n1,
         AddKeyXOR2_XORInst_4_0_n1, AddKeyXOR2_XORInst_4_1_n1,
         AddKeyXOR2_XORInst_4_2_n1, AddKeyXOR2_XORInst_4_3_n1,
         AddKeyXOR2_XORInst_5_0_n1, AddKeyXOR2_XORInst_5_1_n1,
         AddKeyXOR2_XORInst_5_2_n1, AddKeyXOR2_XORInst_5_3_n1,
         AddKeyXOR2_XORInst_6_0_n1, AddKeyXOR2_XORInst_6_1_n1,
         AddKeyXOR2_XORInst_6_2_n1, AddKeyXOR2_XORInst_6_3_n1,
         AddKeyXOR2_XORInst_7_0_n1, AddKeyXOR2_XORInst_7_1_n1,
         AddKeyXOR2_XORInst_7_2_n1, AddKeyXOR2_XORInst_7_3_n1,
         AddKeyXOR2_XORInst_8_0_n1, AddKeyXOR2_XORInst_8_1_n1,
         AddKeyXOR2_XORInst_8_2_n1, AddKeyXOR2_XORInst_8_3_n1,
         AddKeyXOR2_XORInst_9_0_n1, AddKeyXOR2_XORInst_9_1_n1,
         AddKeyXOR2_XORInst_9_2_n1, AddKeyXOR2_XORInst_9_3_n1,
         StateReg_s_current_state_reg_63__QN,
         StateReg_s_current_state_reg_62__QN,
         StateReg_s_current_state_reg_61__QN,
         StateReg_s_current_state_reg_60__QN,
         StateReg_s_current_state_reg_59__QN,
         StateReg_s_current_state_reg_58__QN,
         StateReg_s_current_state_reg_57__QN,
         StateReg_s_current_state_reg_56__QN,
         StateReg_s_current_state_reg_55__QN,
         StateReg_s_current_state_reg_54__QN,
         StateReg_s_current_state_reg_53__QN,
         StateReg_s_current_state_reg_52__QN,
         StateReg_s_current_state_reg_51__QN,
         StateReg_s_current_state_reg_50__QN,
         StateReg_s_current_state_reg_49__QN,
         StateReg_s_current_state_reg_48__QN,
         StateReg_s_current_state_reg_47__QN,
         StateReg_s_current_state_reg_46__QN,
         StateReg_s_current_state_reg_45__QN,
         StateReg_s_current_state_reg_44__QN,
         StateReg_s_current_state_reg_43__QN,
         StateReg_s_current_state_reg_42__QN,
         StateReg_s_current_state_reg_41__QN,
         StateReg_s_current_state_reg_40__QN,
         StateReg_s_current_state_reg_39__QN,
         StateReg_s_current_state_reg_38__QN,
         StateReg_s_current_state_reg_37__QN,
         StateReg_s_current_state_reg_36__QN,
         StateReg_s_current_state_reg_35__QN,
         StateReg_s_current_state_reg_34__QN,
         StateReg_s_current_state_reg_33__QN,
         StateReg_s_current_state_reg_32__QN,
         StateReg_s_current_state_reg_31__QN,
         StateReg_s_current_state_reg_30__QN,
         StateReg_s_current_state_reg_29__QN,
         StateReg_s_current_state_reg_28__QN,
         StateReg_s_current_state_reg_27__QN,
         StateReg_s_current_state_reg_26__QN,
         StateReg_s_current_state_reg_25__QN,
         StateReg_s_current_state_reg_24__QN,
         StateReg_s_current_state_reg_23__QN,
         StateReg_s_current_state_reg_22__QN,
         StateReg_s_current_state_reg_21__QN,
         StateReg_s_current_state_reg_20__QN,
         StateReg_s_current_state_reg_19__QN,
         StateReg_s_current_state_reg_18__QN,
         StateReg_s_current_state_reg_17__QN,
         StateReg_s_current_state_reg_16__QN,
         StateReg_s_current_state_reg_15__QN,
         StateReg_s_current_state_reg_14__QN,
         StateReg_s_current_state_reg_13__QN,
         StateReg_s_current_state_reg_12__QN,
         StateReg_s_current_state_reg_11__QN,
         StateReg_s_current_state_reg_10__QN,
         StateReg_s_current_state_reg_9__QN,
         StateReg_s_current_state_reg_8__QN,
         StateReg_s_current_state_reg_7__QN,
         StateReg_s_current_state_reg_6__QN,
         StateReg_s_current_state_reg_5__QN,
         StateReg_s_current_state_reg_4__QN,
         StateReg_s_current_state_reg_3__QN,
         StateReg_s_current_state_reg_2__QN,
         StateReg_s_current_state_reg_1__QN,
         StateReg_s_current_state_reg_0__QN, SubCellInst_SboxInst_0_n15,
         SubCellInst_SboxInst_0_n14, SubCellInst_SboxInst_0_n13,
         SubCellInst_SboxInst_0_n12, SubCellInst_SboxInst_0_n11,
         SubCellInst_SboxInst_0_n10, SubCellInst_SboxInst_0_n9,
         SubCellInst_SboxInst_0_n8, SubCellInst_SboxInst_0_n7,
         SubCellInst_SboxInst_0_n6, SubCellInst_SboxInst_0_n5,
         SubCellInst_SboxInst_0_n4, SubCellInst_SboxInst_0_n3,
         SubCellInst_SboxInst_0_n2, SubCellInst_SboxInst_0_n1,
         SubCellInst_SboxInst_1_n15, SubCellInst_SboxInst_1_n14,
         SubCellInst_SboxInst_1_n13, SubCellInst_SboxInst_1_n12,
         SubCellInst_SboxInst_1_n11, SubCellInst_SboxInst_1_n10,
         SubCellInst_SboxInst_1_n9, SubCellInst_SboxInst_1_n8,
         SubCellInst_SboxInst_1_n7, SubCellInst_SboxInst_1_n6,
         SubCellInst_SboxInst_1_n5, SubCellInst_SboxInst_1_n4,
         SubCellInst_SboxInst_1_n3, SubCellInst_SboxInst_1_n2,
         SubCellInst_SboxInst_1_n1, SubCellInst_SboxInst_2_n15,
         SubCellInst_SboxInst_2_n14, SubCellInst_SboxInst_2_n13,
         SubCellInst_SboxInst_2_n12, SubCellInst_SboxInst_2_n11,
         SubCellInst_SboxInst_2_n10, SubCellInst_SboxInst_2_n9,
         SubCellInst_SboxInst_2_n8, SubCellInst_SboxInst_2_n7,
         SubCellInst_SboxInst_2_n6, SubCellInst_SboxInst_2_n5,
         SubCellInst_SboxInst_2_n4, SubCellInst_SboxInst_2_n3,
         SubCellInst_SboxInst_2_n2, SubCellInst_SboxInst_2_n1,
         SubCellInst_SboxInst_3_n15, SubCellInst_SboxInst_3_n14,
         SubCellInst_SboxInst_3_n13, SubCellInst_SboxInst_3_n12,
         SubCellInst_SboxInst_3_n11, SubCellInst_SboxInst_3_n10,
         SubCellInst_SboxInst_3_n9, SubCellInst_SboxInst_3_n8,
         SubCellInst_SboxInst_3_n7, SubCellInst_SboxInst_3_n6,
         SubCellInst_SboxInst_3_n5, SubCellInst_SboxInst_3_n4,
         SubCellInst_SboxInst_3_n3, SubCellInst_SboxInst_3_n2,
         SubCellInst_SboxInst_3_n1, SubCellInst_SboxInst_4_n15,
         SubCellInst_SboxInst_4_n14, SubCellInst_SboxInst_4_n13,
         SubCellInst_SboxInst_4_n12, SubCellInst_SboxInst_4_n11,
         SubCellInst_SboxInst_4_n10, SubCellInst_SboxInst_4_n9,
         SubCellInst_SboxInst_4_n8, SubCellInst_SboxInst_4_n7,
         SubCellInst_SboxInst_4_n6, SubCellInst_SboxInst_4_n5,
         SubCellInst_SboxInst_4_n4, SubCellInst_SboxInst_4_n3,
         SubCellInst_SboxInst_4_n2, SubCellInst_SboxInst_4_n1,
         SubCellInst_SboxInst_5_n15, SubCellInst_SboxInst_5_n14,
         SubCellInst_SboxInst_5_n13, SubCellInst_SboxInst_5_n12,
         SubCellInst_SboxInst_5_n11, SubCellInst_SboxInst_5_n10,
         SubCellInst_SboxInst_5_n9, SubCellInst_SboxInst_5_n8,
         SubCellInst_SboxInst_5_n7, SubCellInst_SboxInst_5_n6,
         SubCellInst_SboxInst_5_n5, SubCellInst_SboxInst_5_n4,
         SubCellInst_SboxInst_5_n3, SubCellInst_SboxInst_5_n2,
         SubCellInst_SboxInst_5_n1, SubCellInst_SboxInst_6_n15,
         SubCellInst_SboxInst_6_n14, SubCellInst_SboxInst_6_n13,
         SubCellInst_SboxInst_6_n12, SubCellInst_SboxInst_6_n11,
         SubCellInst_SboxInst_6_n10, SubCellInst_SboxInst_6_n9,
         SubCellInst_SboxInst_6_n8, SubCellInst_SboxInst_6_n7,
         SubCellInst_SboxInst_6_n6, SubCellInst_SboxInst_6_n5,
         SubCellInst_SboxInst_6_n4, SubCellInst_SboxInst_6_n3,
         SubCellInst_SboxInst_6_n2, SubCellInst_SboxInst_6_n1,
         SubCellInst_SboxInst_7_n15, SubCellInst_SboxInst_7_n14,
         SubCellInst_SboxInst_7_n13, SubCellInst_SboxInst_7_n12,
         SubCellInst_SboxInst_7_n11, SubCellInst_SboxInst_7_n10,
         SubCellInst_SboxInst_7_n9, SubCellInst_SboxInst_7_n8,
         SubCellInst_SboxInst_7_n7, SubCellInst_SboxInst_7_n6,
         SubCellInst_SboxInst_7_n5, SubCellInst_SboxInst_7_n4,
         SubCellInst_SboxInst_7_n3, SubCellInst_SboxInst_7_n2,
         SubCellInst_SboxInst_7_n1, SubCellInst_SboxInst_8_n15,
         SubCellInst_SboxInst_8_n14, SubCellInst_SboxInst_8_n13,
         SubCellInst_SboxInst_8_n12, SubCellInst_SboxInst_8_n11,
         SubCellInst_SboxInst_8_n10, SubCellInst_SboxInst_8_n9,
         SubCellInst_SboxInst_8_n8, SubCellInst_SboxInst_8_n7,
         SubCellInst_SboxInst_8_n6, SubCellInst_SboxInst_8_n5,
         SubCellInst_SboxInst_8_n4, SubCellInst_SboxInst_8_n3,
         SubCellInst_SboxInst_8_n2, SubCellInst_SboxInst_8_n1,
         SubCellInst_SboxInst_9_n15, SubCellInst_SboxInst_9_n14,
         SubCellInst_SboxInst_9_n13, SubCellInst_SboxInst_9_n12,
         SubCellInst_SboxInst_9_n11, SubCellInst_SboxInst_9_n10,
         SubCellInst_SboxInst_9_n9, SubCellInst_SboxInst_9_n8,
         SubCellInst_SboxInst_9_n7, SubCellInst_SboxInst_9_n6,
         SubCellInst_SboxInst_9_n5, SubCellInst_SboxInst_9_n4,
         SubCellInst_SboxInst_9_n3, SubCellInst_SboxInst_9_n2,
         SubCellInst_SboxInst_9_n1, SubCellInst_SboxInst_10_n15,
         SubCellInst_SboxInst_10_n14, SubCellInst_SboxInst_10_n13,
         SubCellInst_SboxInst_10_n12, SubCellInst_SboxInst_10_n11,
         SubCellInst_SboxInst_10_n10, SubCellInst_SboxInst_10_n9,
         SubCellInst_SboxInst_10_n8, SubCellInst_SboxInst_10_n7,
         SubCellInst_SboxInst_10_n6, SubCellInst_SboxInst_10_n5,
         SubCellInst_SboxInst_10_n4, SubCellInst_SboxInst_10_n3,
         SubCellInst_SboxInst_10_n2, SubCellInst_SboxInst_10_n1,
         SubCellInst_SboxInst_11_n15, SubCellInst_SboxInst_11_n14,
         SubCellInst_SboxInst_11_n13, SubCellInst_SboxInst_11_n12,
         SubCellInst_SboxInst_11_n11, SubCellInst_SboxInst_11_n10,
         SubCellInst_SboxInst_11_n9, SubCellInst_SboxInst_11_n8,
         SubCellInst_SboxInst_11_n7, SubCellInst_SboxInst_11_n6,
         SubCellInst_SboxInst_11_n5, SubCellInst_SboxInst_11_n4,
         SubCellInst_SboxInst_11_n3, SubCellInst_SboxInst_11_n2,
         SubCellInst_SboxInst_11_n1, SubCellInst_SboxInst_12_n15,
         SubCellInst_SboxInst_12_n14, SubCellInst_SboxInst_12_n13,
         SubCellInst_SboxInst_12_n12, SubCellInst_SboxInst_12_n11,
         SubCellInst_SboxInst_12_n10, SubCellInst_SboxInst_12_n9,
         SubCellInst_SboxInst_12_n8, SubCellInst_SboxInst_12_n7,
         SubCellInst_SboxInst_12_n6, SubCellInst_SboxInst_12_n5,
         SubCellInst_SboxInst_12_n4, SubCellInst_SboxInst_12_n3,
         SubCellInst_SboxInst_12_n2, SubCellInst_SboxInst_12_n1,
         SubCellInst_SboxInst_13_n15, SubCellInst_SboxInst_13_n14,
         SubCellInst_SboxInst_13_n13, SubCellInst_SboxInst_13_n12,
         SubCellInst_SboxInst_13_n11, SubCellInst_SboxInst_13_n10,
         SubCellInst_SboxInst_13_n9, SubCellInst_SboxInst_13_n8,
         SubCellInst_SboxInst_13_n7, SubCellInst_SboxInst_13_n6,
         SubCellInst_SboxInst_13_n5, SubCellInst_SboxInst_13_n4,
         SubCellInst_SboxInst_13_n3, SubCellInst_SboxInst_13_n2,
         SubCellInst_SboxInst_13_n1, SubCellInst_SboxInst_14_n15,
         SubCellInst_SboxInst_14_n14, SubCellInst_SboxInst_14_n13,
         SubCellInst_SboxInst_14_n12, SubCellInst_SboxInst_14_n11,
         SubCellInst_SboxInst_14_n10, SubCellInst_SboxInst_14_n9,
         SubCellInst_SboxInst_14_n8, SubCellInst_SboxInst_14_n7,
         SubCellInst_SboxInst_14_n6, SubCellInst_SboxInst_14_n5,
         SubCellInst_SboxInst_14_n4, SubCellInst_SboxInst_14_n3,
         SubCellInst_SboxInst_14_n2, SubCellInst_SboxInst_14_n1,
         SubCellInst_SboxInst_15_n15, SubCellInst_SboxInst_15_n14,
         SubCellInst_SboxInst_15_n13, SubCellInst_SboxInst_15_n12,
         SubCellInst_SboxInst_15_n11, SubCellInst_SboxInst_15_n10,
         SubCellInst_SboxInst_15_n9, SubCellInst_SboxInst_15_n8,
         SubCellInst_SboxInst_15_n7, SubCellInst_SboxInst_15_n6,
         SubCellInst_SboxInst_15_n5, SubCellInst_SboxInst_15_n4,
         SubCellInst_SboxInst_15_n3, SubCellInst_SboxInst_15_n2,
         SubCellInst_SboxInst_15_n1, KeyMUX_n9, KeyMUX_n8, KeyMUX_n7,
         FSMRegInst_s_current_state_reg_6__QN,
         FSMRegInst_s_current_state_reg_5__QN,
         FSMRegInst_s_current_state_reg_4__QN,
         FSMRegInst_s_current_state_reg_3__QN,
         FSMRegInst_s_current_state_reg_2__QN,
         FSMRegInst_s_current_state_reg_1__QN,
         FSMRegInst_s_current_state_reg_0__QN, FSMSignalsInst_n5,
         FSMSignalsInst_n4, FSMSignalsInst_n3, FSMSignalsInst_n2,
         FSMSignalsInst_n1, selectsUpdateInst_n3,
         selectsRegInst_s_current_state_reg_1__QN,
         selectsRegInst_s_current_state_reg_0__QN, done_reg_QN;
  wire   [63:0] Feedback;
  wire   [63:32] MCInput;
  wire   [63:0] MCOutput;
  wire   [63:0] SelectedKey;
  wire   [63:0] AddRoundKeyOutput;
  wire   [1:0] selects;
  wire   [6:0] FSMReg;
  wire   [6:0] FSMUpdate;
  wire   [1:0] selectsReg;
  wire   [1:0] selectsNext;

  MUX2_X1 InputMUX_MUXInst_0_U1 ( .A(Feedback[0]), .B(plaintext[0]), .S(rst), .Z(
        MCOutput[0]) );
  MUX2_X1 InputMUX_MUXInst_1_U1 ( .A(Feedback[1]), .B(plaintext[1]), .S(rst), .Z(
        MCOutput[1]) );
  MUX2_X1 InputMUX_MUXInst_2_U1 ( .A(Feedback[2]), .B(plaintext[2]), .S(rst), .Z(
        MCOutput[2]) );
  MUX2_X1 InputMUX_MUXInst_3_U1 ( .A(Feedback[3]), .B(plaintext[3]), .S(rst), .Z(
        MCOutput[3]) );
  MUX2_X1 InputMUX_MUXInst_4_U1 ( .A(Feedback[4]), .B(plaintext[4]), .S(rst), .Z(
        MCOutput[4]) );
  MUX2_X1 InputMUX_MUXInst_5_U1 ( .A(Feedback[5]), .B(plaintext[5]), .S(rst), .Z(
        MCOutput[5]) );
  MUX2_X1 InputMUX_MUXInst_6_U1 ( .A(Feedback[6]), .B(plaintext[6]), .S(rst), .Z(
        MCOutput[6]) );
  MUX2_X1 InputMUX_MUXInst_7_U1 ( .A(Feedback[7]), .B(plaintext[7]), .S(rst), .Z(
        MCOutput[7]) );
  MUX2_X1 InputMUX_MUXInst_8_U1 ( .A(Feedback[8]), .B(plaintext[8]), .S(rst), .Z(
        MCOutput[8]) );
  MUX2_X1 InputMUX_MUXInst_9_U1 ( .A(Feedback[9]), .B(plaintext[9]), .S(rst), .Z(
        MCOutput[9]) );
  MUX2_X1 InputMUX_MUXInst_10_U1 ( .A(Feedback[10]), .B(plaintext[10]), .S(rst), 
        .Z(MCOutput[10]) );
  MUX2_X1 InputMUX_MUXInst_11_U1 ( .A(Feedback[11]), .B(plaintext[11]), .S(rst), 
        .Z(MCOutput[11]) );
  MUX2_X1 InputMUX_MUXInst_12_U1 ( .A(Feedback[12]), .B(plaintext[12]), .S(rst), 
        .Z(MCOutput[12]) );
  MUX2_X1 InputMUX_MUXInst_13_U1 ( .A(Feedback[13]), .B(plaintext[13]), .S(rst), 
        .Z(MCOutput[13]) );
  MUX2_X1 InputMUX_MUXInst_14_U1 ( .A(Feedback[14]), .B(plaintext[14]), .S(rst), 
        .Z(MCOutput[14]) );
  MUX2_X1 InputMUX_MUXInst_15_U1 ( .A(Feedback[15]), .B(plaintext[15]), .S(rst), 
        .Z(MCOutput[15]) );
  MUX2_X1 InputMUX_MUXInst_16_U1 ( .A(Feedback[16]), .B(plaintext[16]), .S(rst), 
        .Z(MCOutput[16]) );
  MUX2_X1 InputMUX_MUXInst_17_U1 ( .A(Feedback[17]), .B(plaintext[17]), .S(rst), 
        .Z(MCOutput[17]) );
  MUX2_X1 InputMUX_MUXInst_18_U1 ( .A(Feedback[18]), .B(plaintext[18]), .S(rst), 
        .Z(MCOutput[18]) );
  MUX2_X1 InputMUX_MUXInst_19_U1 ( .A(Feedback[19]), .B(plaintext[19]), .S(rst), 
        .Z(MCOutput[19]) );
  MUX2_X1 InputMUX_MUXInst_20_U1 ( .A(Feedback[20]), .B(plaintext[20]), .S(rst), 
        .Z(MCOutput[20]) );
  MUX2_X1 InputMUX_MUXInst_21_U1 ( .A(Feedback[21]), .B(plaintext[21]), .S(rst), 
        .Z(MCOutput[21]) );
  MUX2_X1 InputMUX_MUXInst_22_U1 ( .A(Feedback[22]), .B(plaintext[22]), .S(rst), 
        .Z(MCOutput[22]) );
  MUX2_X1 InputMUX_MUXInst_23_U1 ( .A(Feedback[23]), .B(plaintext[23]), .S(rst), 
        .Z(MCOutput[23]) );
  MUX2_X1 InputMUX_MUXInst_24_U1 ( .A(Feedback[24]), .B(plaintext[24]), .S(rst), 
        .Z(MCOutput[24]) );
  MUX2_X1 InputMUX_MUXInst_25_U1 ( .A(Feedback[25]), .B(plaintext[25]), .S(rst), 
        .Z(MCOutput[25]) );
  MUX2_X1 InputMUX_MUXInst_26_U1 ( .A(Feedback[26]), .B(plaintext[26]), .S(rst), 
        .Z(MCOutput[26]) );
  MUX2_X1 InputMUX_MUXInst_27_U1 ( .A(Feedback[27]), .B(plaintext[27]), .S(rst), 
        .Z(MCOutput[27]) );
  MUX2_X1 InputMUX_MUXInst_28_U1 ( .A(Feedback[28]), .B(plaintext[28]), .S(rst), 
        .Z(MCOutput[28]) );
  MUX2_X1 InputMUX_MUXInst_29_U1 ( .A(Feedback[29]), .B(plaintext[29]), .S(rst), 
        .Z(MCOutput[29]) );
  MUX2_X1 InputMUX_MUXInst_30_U1 ( .A(Feedback[30]), .B(plaintext[30]), .S(rst), 
        .Z(MCOutput[30]) );
  MUX2_X1 InputMUX_MUXInst_31_U1 ( .A(Feedback[31]), .B(plaintext[31]), .S(rst), 
        .Z(MCOutput[31]) );
  MUX2_X1 InputMUX_MUXInst_32_U1 ( .A(Feedback[32]), .B(plaintext[32]), .S(rst), 
        .Z(MCInput[32]) );
  MUX2_X1 InputMUX_MUXInst_33_U1 ( .A(Feedback[33]), .B(plaintext[33]), .S(rst), 
        .Z(MCInput[33]) );
  MUX2_X1 InputMUX_MUXInst_34_U1 ( .A(Feedback[34]), .B(plaintext[34]), .S(rst), 
        .Z(MCInput[34]) );
  MUX2_X1 InputMUX_MUXInst_35_U1 ( .A(Feedback[35]), .B(plaintext[35]), .S(rst), 
        .Z(MCInput[35]) );
  MUX2_X1 InputMUX_MUXInst_36_U1 ( .A(Feedback[36]), .B(plaintext[36]), .S(rst), 
        .Z(MCInput[36]) );
  MUX2_X1 InputMUX_MUXInst_37_U1 ( .A(Feedback[37]), .B(plaintext[37]), .S(rst), 
        .Z(MCInput[37]) );
  MUX2_X1 InputMUX_MUXInst_38_U1 ( .A(Feedback[38]), .B(plaintext[38]), .S(rst), 
        .Z(MCInput[38]) );
  MUX2_X1 InputMUX_MUXInst_39_U1 ( .A(Feedback[39]), .B(plaintext[39]), .S(rst), 
        .Z(MCInput[39]) );
  MUX2_X1 InputMUX_MUXInst_40_U1 ( .A(Feedback[40]), .B(plaintext[40]), .S(rst), 
        .Z(MCInput[40]) );
  MUX2_X1 InputMUX_MUXInst_41_U1 ( .A(Feedback[41]), .B(plaintext[41]), .S(rst), 
        .Z(MCInput[41]) );
  MUX2_X1 InputMUX_MUXInst_42_U1 ( .A(Feedback[42]), .B(plaintext[42]), .S(rst), 
        .Z(MCInput[42]) );
  MUX2_X1 InputMUX_MUXInst_43_U1 ( .A(Feedback[43]), .B(plaintext[43]), .S(rst), 
        .Z(MCInput[43]) );
  MUX2_X1 InputMUX_MUXInst_44_U1 ( .A(Feedback[44]), .B(plaintext[44]), .S(rst), 
        .Z(MCInput[44]) );
  MUX2_X1 InputMUX_MUXInst_45_U1 ( .A(Feedback[45]), .B(plaintext[45]), .S(rst), 
        .Z(MCInput[45]) );
  MUX2_X1 InputMUX_MUXInst_46_U1 ( .A(Feedback[46]), .B(plaintext[46]), .S(rst), 
        .Z(MCInput[46]) );
  MUX2_X1 InputMUX_MUXInst_47_U1 ( .A(Feedback[47]), .B(plaintext[47]), .S(rst), 
        .Z(MCInput[47]) );
  MUX2_X1 InputMUX_MUXInst_48_U1 ( .A(Feedback[48]), .B(plaintext[48]), .S(rst), 
        .Z(MCInput[48]) );
  MUX2_X1 InputMUX_MUXInst_49_U1 ( .A(Feedback[49]), .B(plaintext[49]), .S(rst), 
        .Z(MCInput[49]) );
  MUX2_X1 InputMUX_MUXInst_50_U1 ( .A(Feedback[50]), .B(plaintext[50]), .S(rst), 
        .Z(MCInput[50]) );
  MUX2_X1 InputMUX_MUXInst_51_U1 ( .A(Feedback[51]), .B(plaintext[51]), .S(rst), 
        .Z(MCInput[51]) );
  MUX2_X1 InputMUX_MUXInst_52_U1 ( .A(Feedback[52]), .B(plaintext[52]), .S(rst), 
        .Z(MCInput[52]) );
  MUX2_X1 InputMUX_MUXInst_53_U1 ( .A(Feedback[53]), .B(plaintext[53]), .S(rst), 
        .Z(MCInput[53]) );
  MUX2_X1 InputMUX_MUXInst_54_U1 ( .A(Feedback[54]), .B(plaintext[54]), .S(rst), 
        .Z(MCInput[54]) );
  MUX2_X1 InputMUX_MUXInst_55_U1 ( .A(Feedback[55]), .B(plaintext[55]), .S(rst), 
        .Z(MCInput[55]) );
  MUX2_X1 InputMUX_MUXInst_56_U1 ( .A(Feedback[56]), .B(plaintext[56]), .S(rst), 
        .Z(MCInput[56]) );
  MUX2_X1 InputMUX_MUXInst_57_U1 ( .A(Feedback[57]), .B(plaintext[57]), .S(rst), 
        .Z(MCInput[57]) );
  MUX2_X1 InputMUX_MUXInst_58_U1 ( .A(Feedback[58]), .B(plaintext[58]), .S(rst), 
        .Z(MCInput[58]) );
  MUX2_X1 InputMUX_MUXInst_59_U1 ( .A(Feedback[59]), .B(plaintext[59]), .S(rst), 
        .Z(MCInput[59]) );
  MUX2_X1 InputMUX_MUXInst_60_U1 ( .A(Feedback[60]), .B(plaintext[60]), .S(rst), 
        .Z(MCInput[60]) );
  MUX2_X1 InputMUX_MUXInst_61_U1 ( .A(Feedback[61]), .B(plaintext[61]), .S(rst), 
        .Z(MCInput[61]) );
  MUX2_X1 InputMUX_MUXInst_62_U1 ( .A(Feedback[62]), .B(plaintext[62]), .S(rst), 
        .Z(MCInput[62]) );
  MUX2_X1 InputMUX_MUXInst_63_U1 ( .A(Feedback[63]), .B(plaintext[63]), .S(rst), 
        .Z(MCInput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U3 ( .A(MCInst_XOR_r0_Inst_0_n2), .B(
        MCInst_XOR_r0_Inst_0_n1), .ZN(MCOutput[48]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_0_U2 ( .A(MCOutput[16]), .B(MCOutput[0]), .ZN(
        MCInst_XOR_r0_Inst_0_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_0_U1 ( .A(1'b0), .B(MCInput[48]), .Z(
        MCInst_XOR_r0_Inst_0_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_0_U2 ( .A(MCInst_XOR_r1_Inst_0_n1), .B(
        MCOutput[0]), .ZN(MCOutput[32]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_0_U1 ( .A(1'b0), .B(MCInput[32]), .ZN(
        MCInst_XOR_r1_Inst_0_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U3 ( .A(MCInst_XOR_r0_Inst_1_n2), .B(
        MCInst_XOR_r0_Inst_1_n1), .ZN(MCOutput[49]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_1_U2 ( .A(MCOutput[17]), .B(MCOutput[1]), .ZN(
        MCInst_XOR_r0_Inst_1_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_1_U1 ( .A(1'b0), .B(MCInput[49]), .Z(
        MCInst_XOR_r0_Inst_1_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_1_U2 ( .A(MCInst_XOR_r1_Inst_1_n1), .B(
        MCOutput[1]), .ZN(MCOutput[33]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_1_U1 ( .A(1'b0), .B(MCInput[33]), .ZN(
        MCInst_XOR_r1_Inst_1_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U3 ( .A(MCInst_XOR_r0_Inst_2_n2), .B(
        MCInst_XOR_r0_Inst_2_n1), .ZN(MCOutput[50]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_2_U2 ( .A(MCOutput[18]), .B(MCOutput[2]), .ZN(
        MCInst_XOR_r0_Inst_2_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_2_U1 ( .A(1'b0), .B(MCInput[50]), .Z(
        MCInst_XOR_r0_Inst_2_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_2_U2 ( .A(MCInst_XOR_r1_Inst_2_n1), .B(
        MCOutput[2]), .ZN(MCOutput[34]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_2_U1 ( .A(1'b0), .B(MCInput[34]), .ZN(
        MCInst_XOR_r1_Inst_2_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U3 ( .A(MCInst_XOR_r0_Inst_3_n2), .B(
        MCInst_XOR_r0_Inst_3_n1), .ZN(MCOutput[51]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_3_U2 ( .A(MCOutput[19]), .B(MCOutput[3]), .ZN(
        MCInst_XOR_r0_Inst_3_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_3_U1 ( .A(1'b0), .B(MCInput[51]), .Z(
        MCInst_XOR_r0_Inst_3_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_3_U2 ( .A(MCInst_XOR_r1_Inst_3_n1), .B(
        MCOutput[3]), .ZN(MCOutput[35]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_3_U1 ( .A(1'b0), .B(MCInput[35]), .ZN(
        MCInst_XOR_r1_Inst_3_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U3 ( .A(MCInst_XOR_r0_Inst_4_n2), .B(
        MCInst_XOR_r0_Inst_4_n1), .ZN(MCOutput[52]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_4_U2 ( .A(MCOutput[20]), .B(MCOutput[4]), .ZN(
        MCInst_XOR_r0_Inst_4_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_4_U1 ( .A(1'b0), .B(MCInput[52]), .Z(
        MCInst_XOR_r0_Inst_4_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_4_U2 ( .A(MCInst_XOR_r1_Inst_4_n1), .B(
        MCOutput[4]), .ZN(MCOutput[36]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_4_U1 ( .A(1'b0), .B(MCInput[36]), .ZN(
        MCInst_XOR_r1_Inst_4_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U3 ( .A(MCInst_XOR_r0_Inst_5_n2), .B(
        MCInst_XOR_r0_Inst_5_n1), .ZN(MCOutput[53]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_5_U2 ( .A(MCOutput[21]), .B(MCOutput[5]), .ZN(
        MCInst_XOR_r0_Inst_5_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_5_U1 ( .A(1'b0), .B(MCInput[53]), .Z(
        MCInst_XOR_r0_Inst_5_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_5_U2 ( .A(MCInst_XOR_r1_Inst_5_n1), .B(
        MCOutput[5]), .ZN(MCOutput[37]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_5_U1 ( .A(1'b0), .B(MCInput[37]), .ZN(
        MCInst_XOR_r1_Inst_5_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U3 ( .A(MCInst_XOR_r0_Inst_6_n2), .B(
        MCInst_XOR_r0_Inst_6_n1), .ZN(MCOutput[54]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_6_U2 ( .A(MCOutput[22]), .B(MCOutput[6]), .ZN(
        MCInst_XOR_r0_Inst_6_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_6_U1 ( .A(1'b0), .B(MCInput[54]), .Z(
        MCInst_XOR_r0_Inst_6_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_6_U2 ( .A(MCInst_XOR_r1_Inst_6_n1), .B(
        MCOutput[6]), .ZN(MCOutput[38]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_6_U1 ( .A(1'b0), .B(MCInput[38]), .ZN(
        MCInst_XOR_r1_Inst_6_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U3 ( .A(MCInst_XOR_r0_Inst_7_n2), .B(
        MCInst_XOR_r0_Inst_7_n1), .ZN(MCOutput[55]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_7_U2 ( .A(MCOutput[23]), .B(MCOutput[7]), .ZN(
        MCInst_XOR_r0_Inst_7_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_7_U1 ( .A(1'b0), .B(MCInput[55]), .Z(
        MCInst_XOR_r0_Inst_7_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_7_U2 ( .A(MCInst_XOR_r1_Inst_7_n1), .B(
        MCOutput[7]), .ZN(MCOutput[39]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_7_U1 ( .A(1'b0), .B(MCInput[39]), .ZN(
        MCInst_XOR_r1_Inst_7_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U3 ( .A(MCInst_XOR_r0_Inst_8_n2), .B(
        MCInst_XOR_r0_Inst_8_n1), .ZN(MCOutput[56]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_8_U2 ( .A(MCOutput[24]), .B(MCOutput[8]), .ZN(
        MCInst_XOR_r0_Inst_8_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_8_U1 ( .A(1'b0), .B(MCInput[56]), .Z(
        MCInst_XOR_r0_Inst_8_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_8_U2 ( .A(MCInst_XOR_r1_Inst_8_n1), .B(
        MCOutput[8]), .ZN(MCOutput[40]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_8_U1 ( .A(1'b0), .B(MCInput[40]), .ZN(
        MCInst_XOR_r1_Inst_8_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U3 ( .A(MCInst_XOR_r0_Inst_9_n2), .B(
        MCInst_XOR_r0_Inst_9_n1), .ZN(MCOutput[57]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_9_U2 ( .A(MCOutput[25]), .B(MCOutput[9]), .ZN(
        MCInst_XOR_r0_Inst_9_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_9_U1 ( .A(1'b0), .B(MCInput[57]), .Z(
        MCInst_XOR_r0_Inst_9_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_9_U2 ( .A(MCInst_XOR_r1_Inst_9_n1), .B(
        MCOutput[9]), .ZN(MCOutput[41]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_9_U1 ( .A(1'b0), .B(MCInput[41]), .ZN(
        MCInst_XOR_r1_Inst_9_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U3 ( .A(MCInst_XOR_r0_Inst_10_n2), .B(
        MCInst_XOR_r0_Inst_10_n1), .ZN(MCOutput[58]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_10_U2 ( .A(MCOutput[26]), .B(MCOutput[10]), .ZN(
        MCInst_XOR_r0_Inst_10_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_10_U1 ( .A(1'b0), .B(MCInput[58]), .Z(
        MCInst_XOR_r0_Inst_10_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_10_U2 ( .A(MCInst_XOR_r1_Inst_10_n1), .B(
        MCOutput[10]), .ZN(MCOutput[42]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_10_U1 ( .A(1'b0), .B(MCInput[42]), .ZN(
        MCInst_XOR_r1_Inst_10_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U3 ( .A(MCInst_XOR_r0_Inst_11_n2), .B(
        MCInst_XOR_r0_Inst_11_n1), .ZN(MCOutput[59]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_11_U2 ( .A(MCOutput[27]), .B(MCOutput[11]), .ZN(
        MCInst_XOR_r0_Inst_11_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_11_U1 ( .A(1'b0), .B(MCInput[59]), .Z(
        MCInst_XOR_r0_Inst_11_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_11_U2 ( .A(MCInst_XOR_r1_Inst_11_n1), .B(
        MCOutput[11]), .ZN(MCOutput[43]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_11_U1 ( .A(1'b0), .B(MCInput[43]), .ZN(
        MCInst_XOR_r1_Inst_11_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U3 ( .A(MCInst_XOR_r0_Inst_12_n2), .B(
        MCInst_XOR_r0_Inst_12_n1), .ZN(MCOutput[60]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_12_U2 ( .A(MCOutput[28]), .B(MCOutput[12]), .ZN(
        MCInst_XOR_r0_Inst_12_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_12_U1 ( .A(1'b0), .B(MCInput[60]), .Z(
        MCInst_XOR_r0_Inst_12_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_12_U2 ( .A(MCInst_XOR_r1_Inst_12_n1), .B(
        MCOutput[12]), .ZN(MCOutput[44]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_12_U1 ( .A(1'b0), .B(MCInput[44]), .ZN(
        MCInst_XOR_r1_Inst_12_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U3 ( .A(MCInst_XOR_r0_Inst_13_n2), .B(
        MCInst_XOR_r0_Inst_13_n1), .ZN(MCOutput[61]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_13_U2 ( .A(MCOutput[29]), .B(MCOutput[13]), .ZN(
        MCInst_XOR_r0_Inst_13_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_13_U1 ( .A(1'b0), .B(MCInput[61]), .Z(
        MCInst_XOR_r0_Inst_13_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_13_U2 ( .A(MCInst_XOR_r1_Inst_13_n1), .B(
        MCOutput[13]), .ZN(MCOutput[45]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_13_U1 ( .A(1'b0), .B(MCInput[45]), .ZN(
        MCInst_XOR_r1_Inst_13_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U3 ( .A(MCInst_XOR_r0_Inst_14_n2), .B(
        MCInst_XOR_r0_Inst_14_n1), .ZN(MCOutput[62]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_14_U2 ( .A(MCOutput[30]), .B(MCOutput[14]), .ZN(
        MCInst_XOR_r0_Inst_14_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_14_U1 ( .A(1'b0), .B(MCInput[62]), .Z(
        MCInst_XOR_r0_Inst_14_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_14_U2 ( .A(MCInst_XOR_r1_Inst_14_n1), .B(
        MCOutput[14]), .ZN(MCOutput[46]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_14_U1 ( .A(1'b0), .B(MCInput[46]), .ZN(
        MCInst_XOR_r1_Inst_14_n1) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U3 ( .A(MCInst_XOR_r0_Inst_15_n2), .B(
        MCInst_XOR_r0_Inst_15_n1), .ZN(MCOutput[63]) );
  XNOR2_X1 MCInst_XOR_r0_Inst_15_U2 ( .A(MCOutput[31]), .B(MCOutput[15]), .ZN(
        MCInst_XOR_r0_Inst_15_n1) );
  XOR2_X1 MCInst_XOR_r0_Inst_15_U1 ( .A(1'b0), .B(MCInput[63]), .Z(
        MCInst_XOR_r0_Inst_15_n2) );
  XNOR2_X1 MCInst_XOR_r1_Inst_15_U2 ( .A(MCInst_XOR_r1_Inst_15_n1), .B(
        MCOutput[15]), .ZN(MCOutput[47]) );
  XNOR2_X1 MCInst_XOR_r1_Inst_15_U1 ( .A(1'b0), .B(MCInput[47]), .ZN(
        MCInst_XOR_r1_Inst_15_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_0_U2 ( .A(AddKeyXOR1_XORInst_0_0_n1), .B(
        SelectedKey[48]), .ZN(AddRoundKeyOutput[48]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[48]), .ZN(
        AddKeyXOR1_XORInst_0_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_1_U2 ( .A(AddKeyXOR1_XORInst_0_1_n1), .B(
        SelectedKey[49]), .ZN(AddRoundKeyOutput[49]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[49]), .ZN(
        AddKeyXOR1_XORInst_0_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_2_U2 ( .A(AddKeyXOR1_XORInst_0_2_n1), .B(
        SelectedKey[50]), .ZN(AddRoundKeyOutput[50]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[50]), .ZN(
        AddKeyXOR1_XORInst_0_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_3_U2 ( .A(AddKeyXOR1_XORInst_0_3_n1), .B(
        SelectedKey[51]), .ZN(AddRoundKeyOutput[51]) );
  XNOR2_X1 AddKeyXOR1_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[51]), .ZN(
        AddKeyXOR1_XORInst_0_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_0_U2 ( .A(AddKeyXOR1_XORInst_1_0_n1), .B(
        SelectedKey[52]), .ZN(AddRoundKeyOutput[52]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[52]), .ZN(
        AddKeyXOR1_XORInst_1_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_1_U2 ( .A(AddKeyXOR1_XORInst_1_1_n1), .B(
        SelectedKey[53]), .ZN(AddRoundKeyOutput[53]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[53]), .ZN(
        AddKeyXOR1_XORInst_1_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_2_U2 ( .A(AddKeyXOR1_XORInst_1_2_n1), .B(
        SelectedKey[54]), .ZN(AddRoundKeyOutput[54]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[54]), .ZN(
        AddKeyXOR1_XORInst_1_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_3_U2 ( .A(AddKeyXOR1_XORInst_1_3_n1), .B(
        SelectedKey[55]), .ZN(AddRoundKeyOutput[55]) );
  XNOR2_X1 AddKeyXOR1_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[55]), .ZN(
        AddKeyXOR1_XORInst_1_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_0_U2 ( .A(AddKeyXOR1_XORInst_2_0_n1), .B(
        SelectedKey[56]), .ZN(AddRoundKeyOutput[56]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[56]), .ZN(
        AddKeyXOR1_XORInst_2_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_1_U2 ( .A(AddKeyXOR1_XORInst_2_1_n1), .B(
        SelectedKey[57]), .ZN(AddRoundKeyOutput[57]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[57]), .ZN(
        AddKeyXOR1_XORInst_2_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_2_U2 ( .A(AddKeyXOR1_XORInst_2_2_n1), .B(
        SelectedKey[58]), .ZN(AddRoundKeyOutput[58]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[58]), .ZN(
        AddKeyXOR1_XORInst_2_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_3_U2 ( .A(AddKeyXOR1_XORInst_2_3_n1), .B(
        SelectedKey[59]), .ZN(AddRoundKeyOutput[59]) );
  XNOR2_X1 AddKeyXOR1_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[59]), .ZN(
        AddKeyXOR1_XORInst_2_3_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_0_U2 ( .A(AddKeyXOR1_XORInst_3_0_n1), .B(
        SelectedKey[60]), .ZN(AddRoundKeyOutput[60]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[60]), .ZN(
        AddKeyXOR1_XORInst_3_0_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_1_U2 ( .A(AddKeyXOR1_XORInst_3_1_n1), .B(
        SelectedKey[61]), .ZN(AddRoundKeyOutput[61]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[61]), .ZN(
        AddKeyXOR1_XORInst_3_1_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_2_U2 ( .A(AddKeyXOR1_XORInst_3_2_n1), .B(
        SelectedKey[62]), .ZN(AddRoundKeyOutput[62]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[62]), .ZN(
        AddKeyXOR1_XORInst_3_2_n1) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_3_U2 ( .A(AddKeyXOR1_XORInst_3_3_n1), .B(
        SelectedKey[63]), .ZN(AddRoundKeyOutput[63]) );
  XNOR2_X1 AddKeyXOR1_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[63]), .ZN(
        AddKeyXOR1_XORInst_3_3_n1) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U3 ( .A(AddKeyConstXOR_XORInst_0_0_n2), 
        .B(AddKeyConstXOR_XORInst_0_0_n1), .ZN(AddRoundKeyOutput[40]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_0_U2 ( .A(SelectedKey[40]), .B(
        RoundConstant_0), .ZN(AddKeyConstXOR_XORInst_0_0_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[40]), .Z(
        AddKeyConstXOR_XORInst_0_0_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U3 ( .A(AddKeyConstXOR_XORInst_0_1_n2), 
        .B(AddKeyConstXOR_XORInst_0_1_n1), .ZN(AddRoundKeyOutput[41]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_1_U2 ( .A(SelectedKey[41]), .B(
        FSMUpdate[0]), .ZN(AddKeyConstXOR_XORInst_0_1_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[41]), .Z(
        AddKeyConstXOR_XORInst_0_1_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U3 ( .A(AddKeyConstXOR_XORInst_0_2_n2), 
        .B(AddKeyConstXOR_XORInst_0_2_n1), .ZN(AddRoundKeyOutput[42]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_2_U2 ( .A(SelectedKey[42]), .B(
        FSMUpdate[1]), .ZN(AddKeyConstXOR_XORInst_0_2_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[42]), .Z(
        AddKeyConstXOR_XORInst_0_2_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_3_U3 ( .A(AddKeyConstXOR_XORInst_0_3_n2), 
        .B(AddKeyConstXOR_XORInst_0_3_n1), .ZN(AddRoundKeyOutput[43]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_0_3_U2 ( .A(SelectedKey[43]), .B(1'b0), .ZN(
        AddKeyConstXOR_XORInst_0_3_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[43]), .Z(
        AddKeyConstXOR_XORInst_0_3_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U3 ( .A(AddKeyConstXOR_XORInst_1_0_n2), 
        .B(AddKeyConstXOR_XORInst_1_0_n1), .ZN(AddRoundKeyOutput[44]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_0_U2 ( .A(SelectedKey[44]), .B(
        RoundConstant_4_), .ZN(AddKeyConstXOR_XORInst_1_0_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[44]), .Z(
        AddKeyConstXOR_XORInst_1_0_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U3 ( .A(AddKeyConstXOR_XORInst_1_1_n2), 
        .B(AddKeyConstXOR_XORInst_1_1_n1), .ZN(AddRoundKeyOutput[45]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_1_U2 ( .A(SelectedKey[45]), .B(
        FSMUpdate[3]), .ZN(AddKeyConstXOR_XORInst_1_1_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[45]), .Z(
        AddKeyConstXOR_XORInst_1_1_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U3 ( .A(AddKeyConstXOR_XORInst_1_2_n2), 
        .B(AddKeyConstXOR_XORInst_1_2_n1), .ZN(AddRoundKeyOutput[46]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_2_U2 ( .A(SelectedKey[46]), .B(
        FSMUpdate[4]), .ZN(AddKeyConstXOR_XORInst_1_2_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[46]), .Z(
        AddKeyConstXOR_XORInst_1_2_n2) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U3 ( .A(AddKeyConstXOR_XORInst_1_3_n2), 
        .B(AddKeyConstXOR_XORInst_1_3_n1), .ZN(AddRoundKeyOutput[47]) );
  XNOR2_X1 AddKeyConstXOR_XORInst_1_3_U2 ( .A(SelectedKey[47]), .B(
        FSMUpdate[5]), .ZN(AddKeyConstXOR_XORInst_1_3_n1) );
  XOR2_X1 AddKeyConstXOR_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[47]), .Z(
        AddKeyConstXOR_XORInst_1_3_n2) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_0_U2 ( .A(AddKeyXOR2_XORInst_0_0_n1), .B(
        SelectedKey[0]), .ZN(AddRoundKeyOutput[0]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_0_U1 ( .A(1'b0), .B(MCOutput[0]), .ZN(
        AddKeyXOR2_XORInst_0_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_1_U2 ( .A(AddKeyXOR2_XORInst_0_1_n1), .B(
        SelectedKey[1]), .ZN(AddRoundKeyOutput[1]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_1_U1 ( .A(1'b0), .B(MCOutput[1]), .ZN(
        AddKeyXOR2_XORInst_0_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_2_U2 ( .A(AddKeyXOR2_XORInst_0_2_n1), .B(
        SelectedKey[2]), .ZN(AddRoundKeyOutput[2]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_2_U1 ( .A(1'b0), .B(MCOutput[2]), .ZN(
        AddKeyXOR2_XORInst_0_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_3_U2 ( .A(AddKeyXOR2_XORInst_0_3_n1), .B(
        SelectedKey[3]), .ZN(AddRoundKeyOutput[3]) );
  XNOR2_X1 AddKeyXOR2_XORInst_0_3_U1 ( .A(1'b0), .B(MCOutput[3]), .ZN(
        AddKeyXOR2_XORInst_0_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_0_U2 ( .A(AddKeyXOR2_XORInst_1_0_n1), .B(
        SelectedKey[4]), .ZN(AddRoundKeyOutput[4]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_0_U1 ( .A(1'b0), .B(MCOutput[4]), .ZN(
        AddKeyXOR2_XORInst_1_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_1_U2 ( .A(AddKeyXOR2_XORInst_1_1_n1), .B(
        SelectedKey[5]), .ZN(AddRoundKeyOutput[5]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_1_U1 ( .A(1'b0), .B(MCOutput[5]), .ZN(
        AddKeyXOR2_XORInst_1_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_2_U2 ( .A(AddKeyXOR2_XORInst_1_2_n1), .B(
        SelectedKey[6]), .ZN(AddRoundKeyOutput[6]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_2_U1 ( .A(1'b0), .B(MCOutput[6]), .ZN(
        AddKeyXOR2_XORInst_1_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_3_U2 ( .A(AddKeyXOR2_XORInst_1_3_n1), .B(
        SelectedKey[7]), .ZN(AddRoundKeyOutput[7]) );
  XNOR2_X1 AddKeyXOR2_XORInst_1_3_U1 ( .A(1'b0), .B(MCOutput[7]), .ZN(
        AddKeyXOR2_XORInst_1_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_0_U2 ( .A(AddKeyXOR2_XORInst_2_0_n1), .B(
        SelectedKey[8]), .ZN(AddRoundKeyOutput[8]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_0_U1 ( .A(1'b0), .B(MCOutput[8]), .ZN(
        AddKeyXOR2_XORInst_2_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_1_U2 ( .A(AddKeyXOR2_XORInst_2_1_n1), .B(
        SelectedKey[9]), .ZN(AddRoundKeyOutput[9]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_1_U1 ( .A(1'b0), .B(MCOutput[9]), .ZN(
        AddKeyXOR2_XORInst_2_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_2_U2 ( .A(AddKeyXOR2_XORInst_2_2_n1), .B(
        SelectedKey[10]), .ZN(AddRoundKeyOutput[10]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_2_U1 ( .A(1'b0), .B(MCOutput[10]), .ZN(
        AddKeyXOR2_XORInst_2_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_3_U2 ( .A(AddKeyXOR2_XORInst_2_3_n1), .B(
        SelectedKey[11]), .ZN(AddRoundKeyOutput[11]) );
  XNOR2_X1 AddKeyXOR2_XORInst_2_3_U1 ( .A(1'b0), .B(MCOutput[11]), .ZN(
        AddKeyXOR2_XORInst_2_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_0_U2 ( .A(AddKeyXOR2_XORInst_3_0_n1), .B(
        SelectedKey[12]), .ZN(AddRoundKeyOutput[12]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_0_U1 ( .A(1'b0), .B(MCOutput[12]), .ZN(
        AddKeyXOR2_XORInst_3_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_1_U2 ( .A(AddKeyXOR2_XORInst_3_1_n1), .B(
        SelectedKey[13]), .ZN(AddRoundKeyOutput[13]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_1_U1 ( .A(1'b0), .B(MCOutput[13]), .ZN(
        AddKeyXOR2_XORInst_3_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_2_U2 ( .A(AddKeyXOR2_XORInst_3_2_n1), .B(
        SelectedKey[14]), .ZN(AddRoundKeyOutput[14]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_2_U1 ( .A(1'b0), .B(MCOutput[14]), .ZN(
        AddKeyXOR2_XORInst_3_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_3_U2 ( .A(AddKeyXOR2_XORInst_3_3_n1), .B(
        SelectedKey[15]), .ZN(AddRoundKeyOutput[15]) );
  XNOR2_X1 AddKeyXOR2_XORInst_3_3_U1 ( .A(1'b0), .B(MCOutput[15]), .ZN(
        AddKeyXOR2_XORInst_3_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_0_U2 ( .A(AddKeyXOR2_XORInst_4_0_n1), .B(
        SelectedKey[16]), .ZN(AddRoundKeyOutput[16]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_0_U1 ( .A(1'b0), .B(MCOutput[16]), .ZN(
        AddKeyXOR2_XORInst_4_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_1_U2 ( .A(AddKeyXOR2_XORInst_4_1_n1), .B(
        SelectedKey[17]), .ZN(AddRoundKeyOutput[17]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_1_U1 ( .A(1'b0), .B(MCOutput[17]), .ZN(
        AddKeyXOR2_XORInst_4_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_2_U2 ( .A(AddKeyXOR2_XORInst_4_2_n1), .B(
        SelectedKey[18]), .ZN(AddRoundKeyOutput[18]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_2_U1 ( .A(1'b0), .B(MCOutput[18]), .ZN(
        AddKeyXOR2_XORInst_4_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_3_U2 ( .A(AddKeyXOR2_XORInst_4_3_n1), .B(
        SelectedKey[19]), .ZN(AddRoundKeyOutput[19]) );
  XNOR2_X1 AddKeyXOR2_XORInst_4_3_U1 ( .A(1'b0), .B(MCOutput[19]), .ZN(
        AddKeyXOR2_XORInst_4_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_0_U2 ( .A(AddKeyXOR2_XORInst_5_0_n1), .B(
        SelectedKey[20]), .ZN(AddRoundKeyOutput[20]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_0_U1 ( .A(1'b0), .B(MCOutput[20]), .ZN(
        AddKeyXOR2_XORInst_5_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_1_U2 ( .A(AddKeyXOR2_XORInst_5_1_n1), .B(
        SelectedKey[21]), .ZN(AddRoundKeyOutput[21]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_1_U1 ( .A(1'b0), .B(MCOutput[21]), .ZN(
        AddKeyXOR2_XORInst_5_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_2_U2 ( .A(AddKeyXOR2_XORInst_5_2_n1), .B(
        SelectedKey[22]), .ZN(AddRoundKeyOutput[22]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_2_U1 ( .A(1'b0), .B(MCOutput[22]), .ZN(
        AddKeyXOR2_XORInst_5_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_3_U2 ( .A(AddKeyXOR2_XORInst_5_3_n1), .B(
        SelectedKey[23]), .ZN(AddRoundKeyOutput[23]) );
  XNOR2_X1 AddKeyXOR2_XORInst_5_3_U1 ( .A(1'b0), .B(MCOutput[23]), .ZN(
        AddKeyXOR2_XORInst_5_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_0_U2 ( .A(AddKeyXOR2_XORInst_6_0_n1), .B(
        SelectedKey[24]), .ZN(AddRoundKeyOutput[24]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_0_U1 ( .A(1'b0), .B(MCOutput[24]), .ZN(
        AddKeyXOR2_XORInst_6_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_1_U2 ( .A(AddKeyXOR2_XORInst_6_1_n1), .B(
        SelectedKey[25]), .ZN(AddRoundKeyOutput[25]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_1_U1 ( .A(1'b0), .B(MCOutput[25]), .ZN(
        AddKeyXOR2_XORInst_6_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_2_U2 ( .A(AddKeyXOR2_XORInst_6_2_n1), .B(
        SelectedKey[26]), .ZN(AddRoundKeyOutput[26]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_2_U1 ( .A(1'b0), .B(MCOutput[26]), .ZN(
        AddKeyXOR2_XORInst_6_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_3_U2 ( .A(AddKeyXOR2_XORInst_6_3_n1), .B(
        SelectedKey[27]), .ZN(AddRoundKeyOutput[27]) );
  XNOR2_X1 AddKeyXOR2_XORInst_6_3_U1 ( .A(1'b0), .B(MCOutput[27]), .ZN(
        AddKeyXOR2_XORInst_6_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_0_U2 ( .A(AddKeyXOR2_XORInst_7_0_n1), .B(
        SelectedKey[28]), .ZN(AddRoundKeyOutput[28]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_0_U1 ( .A(1'b0), .B(MCOutput[28]), .ZN(
        AddKeyXOR2_XORInst_7_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_1_U2 ( .A(AddKeyXOR2_XORInst_7_1_n1), .B(
        SelectedKey[29]), .ZN(AddRoundKeyOutput[29]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_1_U1 ( .A(1'b0), .B(MCOutput[29]), .ZN(
        AddKeyXOR2_XORInst_7_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_2_U2 ( .A(AddKeyXOR2_XORInst_7_2_n1), .B(
        SelectedKey[30]), .ZN(AddRoundKeyOutput[30]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_2_U1 ( .A(1'b0), .B(MCOutput[30]), .ZN(
        AddKeyXOR2_XORInst_7_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_3_U2 ( .A(AddKeyXOR2_XORInst_7_3_n1), .B(
        SelectedKey[31]), .ZN(AddRoundKeyOutput[31]) );
  XNOR2_X1 AddKeyXOR2_XORInst_7_3_U1 ( .A(1'b0), .B(MCOutput[31]), .ZN(
        AddKeyXOR2_XORInst_7_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_0_U2 ( .A(AddKeyXOR2_XORInst_8_0_n1), .B(
        SelectedKey[32]), .ZN(AddRoundKeyOutput[32]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_0_U1 ( .A(1'b0), .B(MCOutput[32]), .ZN(
        AddKeyXOR2_XORInst_8_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_1_U2 ( .A(AddKeyXOR2_XORInst_8_1_n1), .B(
        SelectedKey[33]), .ZN(AddRoundKeyOutput[33]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_1_U1 ( .A(1'b0), .B(MCOutput[33]), .ZN(
        AddKeyXOR2_XORInst_8_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_2_U2 ( .A(AddKeyXOR2_XORInst_8_2_n1), .B(
        SelectedKey[34]), .ZN(AddRoundKeyOutput[34]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_2_U1 ( .A(1'b0), .B(MCOutput[34]), .ZN(
        AddKeyXOR2_XORInst_8_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_3_U2 ( .A(AddKeyXOR2_XORInst_8_3_n1), .B(
        SelectedKey[35]), .ZN(AddRoundKeyOutput[35]) );
  XNOR2_X1 AddKeyXOR2_XORInst_8_3_U1 ( .A(1'b0), .B(MCOutput[35]), .ZN(
        AddKeyXOR2_XORInst_8_3_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_0_U2 ( .A(AddKeyXOR2_XORInst_9_0_n1), .B(
        SelectedKey[36]), .ZN(AddRoundKeyOutput[36]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_0_U1 ( .A(1'b0), .B(MCOutput[36]), .ZN(
        AddKeyXOR2_XORInst_9_0_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_1_U2 ( .A(AddKeyXOR2_XORInst_9_1_n1), .B(
        SelectedKey[37]), .ZN(AddRoundKeyOutput[37]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_1_U1 ( .A(1'b0), .B(MCOutput[37]), .ZN(
        AddKeyXOR2_XORInst_9_1_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_2_U2 ( .A(AddKeyXOR2_XORInst_9_2_n1), .B(
        SelectedKey[38]), .ZN(AddRoundKeyOutput[38]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_2_U1 ( .A(1'b0), .B(MCOutput[38]), .ZN(
        AddKeyXOR2_XORInst_9_2_n1) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_3_U2 ( .A(AddKeyXOR2_XORInst_9_3_n1), .B(
        SelectedKey[39]), .ZN(AddRoundKeyOutput[39]) );
  XNOR2_X1 AddKeyXOR2_XORInst_9_3_U1 ( .A(1'b0), .B(MCOutput[39]), .ZN(
        AddKeyXOR2_XORInst_9_3_n1) );
  INV_X1 StateReg_s_current_state_reg_63__U1 ( .A(ciphertext[63]), .ZN(
        StateReg_s_current_state_reg_63__QN) );
  DFF_X1 StateReg_s_current_state_reg_63__FF_FF ( .D(AddRoundKeyOutput[63]), 
        .CK(clk), .Q(ciphertext[63]), .QN() );
  INV_X1 StateReg_s_current_state_reg_62__U1 ( .A(ciphertext[62]), .ZN(
        StateReg_s_current_state_reg_62__QN) );
  DFF_X1 StateReg_s_current_state_reg_62__FF_FF ( .D(AddRoundKeyOutput[62]), 
        .CK(clk), .Q(ciphertext[62]), .QN() );
  INV_X1 StateReg_s_current_state_reg_61__U1 ( .A(ciphertext[61]), .ZN(
        StateReg_s_current_state_reg_61__QN) );
  DFF_X1 StateReg_s_current_state_reg_61__FF_FF ( .D(AddRoundKeyOutput[61]), 
        .CK(clk), .Q(ciphertext[61]), .QN() );
  INV_X1 StateReg_s_current_state_reg_60__U1 ( .A(ciphertext[60]), .ZN(
        StateReg_s_current_state_reg_60__QN) );
  DFF_X1 StateReg_s_current_state_reg_60__FF_FF ( .D(AddRoundKeyOutput[60]), 
        .CK(clk), .Q(ciphertext[60]), .QN() );
  INV_X1 StateReg_s_current_state_reg_59__U1 ( .A(ciphertext[59]), .ZN(
        StateReg_s_current_state_reg_59__QN) );
  DFF_X1 StateReg_s_current_state_reg_59__FF_FF ( .D(AddRoundKeyOutput[59]), 
        .CK(clk), .Q(ciphertext[59]), .QN() );
  INV_X1 StateReg_s_current_state_reg_58__U1 ( .A(ciphertext[58]), .ZN(
        StateReg_s_current_state_reg_58__QN) );
  DFF_X1 StateReg_s_current_state_reg_58__FF_FF ( .D(AddRoundKeyOutput[58]), 
        .CK(clk), .Q(ciphertext[58]), .QN() );
  INV_X1 StateReg_s_current_state_reg_57__U1 ( .A(ciphertext[57]), .ZN(
        StateReg_s_current_state_reg_57__QN) );
  DFF_X1 StateReg_s_current_state_reg_57__FF_FF ( .D(AddRoundKeyOutput[57]), 
        .CK(clk), .Q(ciphertext[57]), .QN() );
  INV_X1 StateReg_s_current_state_reg_56__U1 ( .A(ciphertext[56]), .ZN(
        StateReg_s_current_state_reg_56__QN) );
  DFF_X1 StateReg_s_current_state_reg_56__FF_FF ( .D(AddRoundKeyOutput[56]), 
        .CK(clk), .Q(ciphertext[56]), .QN() );
  INV_X1 StateReg_s_current_state_reg_55__U1 ( .A(ciphertext[55]), .ZN(
        StateReg_s_current_state_reg_55__QN) );
  DFF_X1 StateReg_s_current_state_reg_55__FF_FF ( .D(AddRoundKeyOutput[55]), 
        .CK(clk), .Q(ciphertext[55]), .QN() );
  INV_X1 StateReg_s_current_state_reg_54__U1 ( .A(ciphertext[54]), .ZN(
        StateReg_s_current_state_reg_54__QN) );
  DFF_X1 StateReg_s_current_state_reg_54__FF_FF ( .D(AddRoundKeyOutput[54]), 
        .CK(clk), .Q(ciphertext[54]), .QN() );
  INV_X1 StateReg_s_current_state_reg_53__U1 ( .A(ciphertext[53]), .ZN(
        StateReg_s_current_state_reg_53__QN) );
  DFF_X1 StateReg_s_current_state_reg_53__FF_FF ( .D(AddRoundKeyOutput[53]), 
        .CK(clk), .Q(ciphertext[53]), .QN() );
  INV_X1 StateReg_s_current_state_reg_52__U1 ( .A(ciphertext[52]), .ZN(
        StateReg_s_current_state_reg_52__QN) );
  DFF_X1 StateReg_s_current_state_reg_52__FF_FF ( .D(AddRoundKeyOutput[52]), 
        .CK(clk), .Q(ciphertext[52]), .QN() );
  INV_X1 StateReg_s_current_state_reg_51__U1 ( .A(ciphertext[51]), .ZN(
        StateReg_s_current_state_reg_51__QN) );
  DFF_X1 StateReg_s_current_state_reg_51__FF_FF ( .D(AddRoundKeyOutput[51]), 
        .CK(clk), .Q(ciphertext[51]), .QN() );
  INV_X1 StateReg_s_current_state_reg_50__U1 ( .A(ciphertext[50]), .ZN(
        StateReg_s_current_state_reg_50__QN) );
  DFF_X1 StateReg_s_current_state_reg_50__FF_FF ( .D(AddRoundKeyOutput[50]), 
        .CK(clk), .Q(ciphertext[50]), .QN() );
  INV_X1 StateReg_s_current_state_reg_49__U1 ( .A(ciphertext[49]), .ZN(
        StateReg_s_current_state_reg_49__QN) );
  DFF_X1 StateReg_s_current_state_reg_49__FF_FF ( .D(AddRoundKeyOutput[49]), 
        .CK(clk), .Q(ciphertext[49]), .QN() );
  INV_X1 StateReg_s_current_state_reg_48__U1 ( .A(ciphertext[48]), .ZN(
        StateReg_s_current_state_reg_48__QN) );
  DFF_X1 StateReg_s_current_state_reg_48__FF_FF ( .D(AddRoundKeyOutput[48]), 
        .CK(clk), .Q(ciphertext[48]), .QN() );
  INV_X1 StateReg_s_current_state_reg_47__U1 ( .A(ciphertext[47]), .ZN(
        StateReg_s_current_state_reg_47__QN) );
  DFF_X1 StateReg_s_current_state_reg_47__FF_FF ( .D(AddRoundKeyOutput[47]), 
        .CK(clk), .Q(ciphertext[47]), .QN() );
  INV_X1 StateReg_s_current_state_reg_46__U1 ( .A(ciphertext[46]), .ZN(
        StateReg_s_current_state_reg_46__QN) );
  DFF_X1 StateReg_s_current_state_reg_46__FF_FF ( .D(AddRoundKeyOutput[46]), 
        .CK(clk), .Q(ciphertext[46]), .QN() );
  INV_X1 StateReg_s_current_state_reg_45__U1 ( .A(ciphertext[45]), .ZN(
        StateReg_s_current_state_reg_45__QN) );
  DFF_X1 StateReg_s_current_state_reg_45__FF_FF ( .D(AddRoundKeyOutput[45]), 
        .CK(clk), .Q(ciphertext[45]), .QN() );
  INV_X1 StateReg_s_current_state_reg_44__U1 ( .A(ciphertext[44]), .ZN(
        StateReg_s_current_state_reg_44__QN) );
  DFF_X1 StateReg_s_current_state_reg_44__FF_FF ( .D(AddRoundKeyOutput[44]), 
        .CK(clk), .Q(ciphertext[44]), .QN() );
  INV_X1 StateReg_s_current_state_reg_43__U1 ( .A(ciphertext[43]), .ZN(
        StateReg_s_current_state_reg_43__QN) );
  DFF_X1 StateReg_s_current_state_reg_43__FF_FF ( .D(AddRoundKeyOutput[43]), 
        .CK(clk), .Q(ciphertext[43]), .QN() );
  INV_X1 StateReg_s_current_state_reg_42__U1 ( .A(ciphertext[42]), .ZN(
        StateReg_s_current_state_reg_42__QN) );
  DFF_X1 StateReg_s_current_state_reg_42__FF_FF ( .D(AddRoundKeyOutput[42]), 
        .CK(clk), .Q(ciphertext[42]), .QN() );
  INV_X1 StateReg_s_current_state_reg_41__U1 ( .A(ciphertext[41]), .ZN(
        StateReg_s_current_state_reg_41__QN) );
  DFF_X1 StateReg_s_current_state_reg_41__FF_FF ( .D(AddRoundKeyOutput[41]), 
        .CK(clk), .Q(ciphertext[41]), .QN() );
  INV_X1 StateReg_s_current_state_reg_40__U1 ( .A(ciphertext[40]), .ZN(
        StateReg_s_current_state_reg_40__QN) );
  DFF_X1 StateReg_s_current_state_reg_40__FF_FF ( .D(AddRoundKeyOutput[40]), 
        .CK(clk), .Q(ciphertext[40]), .QN() );
  INV_X1 StateReg_s_current_state_reg_39__U1 ( .A(ciphertext[39]), .ZN(
        StateReg_s_current_state_reg_39__QN) );
  DFF_X1 StateReg_s_current_state_reg_39__FF_FF ( .D(AddRoundKeyOutput[39]), 
        .CK(clk), .Q(ciphertext[39]), .QN() );
  INV_X1 StateReg_s_current_state_reg_38__U1 ( .A(ciphertext[38]), .ZN(
        StateReg_s_current_state_reg_38__QN) );
  DFF_X1 StateReg_s_current_state_reg_38__FF_FF ( .D(AddRoundKeyOutput[38]), 
        .CK(clk), .Q(ciphertext[38]), .QN() );
  INV_X1 StateReg_s_current_state_reg_37__U1 ( .A(ciphertext[37]), .ZN(
        StateReg_s_current_state_reg_37__QN) );
  DFF_X1 StateReg_s_current_state_reg_37__FF_FF ( .D(AddRoundKeyOutput[37]), 
        .CK(clk), .Q(ciphertext[37]), .QN() );
  INV_X1 StateReg_s_current_state_reg_36__U1 ( .A(ciphertext[36]), .ZN(
        StateReg_s_current_state_reg_36__QN) );
  DFF_X1 StateReg_s_current_state_reg_36__FF_FF ( .D(AddRoundKeyOutput[36]), 
        .CK(clk), .Q(ciphertext[36]), .QN() );
  INV_X1 StateReg_s_current_state_reg_35__U1 ( .A(ciphertext[35]), .ZN(
        StateReg_s_current_state_reg_35__QN) );
  DFF_X1 StateReg_s_current_state_reg_35__FF_FF ( .D(AddRoundKeyOutput[35]), 
        .CK(clk), .Q(ciphertext[35]), .QN() );
  INV_X1 StateReg_s_current_state_reg_34__U1 ( .A(ciphertext[34]), .ZN(
        StateReg_s_current_state_reg_34__QN) );
  DFF_X1 StateReg_s_current_state_reg_34__FF_FF ( .D(AddRoundKeyOutput[34]), 
        .CK(clk), .Q(ciphertext[34]), .QN() );
  INV_X1 StateReg_s_current_state_reg_33__U1 ( .A(ciphertext[33]), .ZN(
        StateReg_s_current_state_reg_33__QN) );
  DFF_X1 StateReg_s_current_state_reg_33__FF_FF ( .D(AddRoundKeyOutput[33]), 
        .CK(clk), .Q(ciphertext[33]), .QN() );
  INV_X1 StateReg_s_current_state_reg_32__U1 ( .A(ciphertext[32]), .ZN(
        StateReg_s_current_state_reg_32__QN) );
  DFF_X1 StateReg_s_current_state_reg_32__FF_FF ( .D(AddRoundKeyOutput[32]), 
        .CK(clk), .Q(ciphertext[32]), .QN() );
  INV_X1 StateReg_s_current_state_reg_31__U1 ( .A(ciphertext[31]), .ZN(
        StateReg_s_current_state_reg_31__QN) );
  DFF_X1 StateReg_s_current_state_reg_31__FF_FF ( .D(AddRoundKeyOutput[31]), 
        .CK(clk), .Q(ciphertext[31]), .QN() );
  INV_X1 StateReg_s_current_state_reg_30__U1 ( .A(ciphertext[30]), .ZN(
        StateReg_s_current_state_reg_30__QN) );
  DFF_X1 StateReg_s_current_state_reg_30__FF_FF ( .D(AddRoundKeyOutput[30]), 
        .CK(clk), .Q(ciphertext[30]), .QN() );
  INV_X1 StateReg_s_current_state_reg_29__U1 ( .A(ciphertext[29]), .ZN(
        StateReg_s_current_state_reg_29__QN) );
  DFF_X1 StateReg_s_current_state_reg_29__FF_FF ( .D(AddRoundKeyOutput[29]), 
        .CK(clk), .Q(ciphertext[29]), .QN() );
  INV_X1 StateReg_s_current_state_reg_28__U1 ( .A(ciphertext[28]), .ZN(
        StateReg_s_current_state_reg_28__QN) );
  DFF_X1 StateReg_s_current_state_reg_28__FF_FF ( .D(AddRoundKeyOutput[28]), 
        .CK(clk), .Q(ciphertext[28]), .QN() );
  INV_X1 StateReg_s_current_state_reg_27__U1 ( .A(ciphertext[27]), .ZN(
        StateReg_s_current_state_reg_27__QN) );
  DFF_X1 StateReg_s_current_state_reg_27__FF_FF ( .D(AddRoundKeyOutput[27]), 
        .CK(clk), .Q(ciphertext[27]), .QN() );
  INV_X1 StateReg_s_current_state_reg_26__U1 ( .A(ciphertext[26]), .ZN(
        StateReg_s_current_state_reg_26__QN) );
  DFF_X1 StateReg_s_current_state_reg_26__FF_FF ( .D(AddRoundKeyOutput[26]), 
        .CK(clk), .Q(ciphertext[26]), .QN() );
  INV_X1 StateReg_s_current_state_reg_25__U1 ( .A(ciphertext[25]), .ZN(
        StateReg_s_current_state_reg_25__QN) );
  DFF_X1 StateReg_s_current_state_reg_25__FF_FF ( .D(AddRoundKeyOutput[25]), 
        .CK(clk), .Q(ciphertext[25]), .QN() );
  INV_X1 StateReg_s_current_state_reg_24__U1 ( .A(ciphertext[24]), .ZN(
        StateReg_s_current_state_reg_24__QN) );
  DFF_X1 StateReg_s_current_state_reg_24__FF_FF ( .D(AddRoundKeyOutput[24]), 
        .CK(clk), .Q(ciphertext[24]), .QN() );
  INV_X1 StateReg_s_current_state_reg_23__U1 ( .A(ciphertext[23]), .ZN(
        StateReg_s_current_state_reg_23__QN) );
  DFF_X1 StateReg_s_current_state_reg_23__FF_FF ( .D(AddRoundKeyOutput[23]), 
        .CK(clk), .Q(ciphertext[23]), .QN() );
  INV_X1 StateReg_s_current_state_reg_22__U1 ( .A(ciphertext[22]), .ZN(
        StateReg_s_current_state_reg_22__QN) );
  DFF_X1 StateReg_s_current_state_reg_22__FF_FF ( .D(AddRoundKeyOutput[22]), 
        .CK(clk), .Q(ciphertext[22]), .QN() );
  INV_X1 StateReg_s_current_state_reg_21__U1 ( .A(ciphertext[21]), .ZN(
        StateReg_s_current_state_reg_21__QN) );
  DFF_X1 StateReg_s_current_state_reg_21__FF_FF ( .D(AddRoundKeyOutput[21]), 
        .CK(clk), .Q(ciphertext[21]), .QN() );
  INV_X1 StateReg_s_current_state_reg_20__U1 ( .A(ciphertext[20]), .ZN(
        StateReg_s_current_state_reg_20__QN) );
  DFF_X1 StateReg_s_current_state_reg_20__FF_FF ( .D(AddRoundKeyOutput[20]), 
        .CK(clk), .Q(ciphertext[20]), .QN() );
  INV_X1 StateReg_s_current_state_reg_19__U1 ( .A(ciphertext[19]), .ZN(
        StateReg_s_current_state_reg_19__QN) );
  DFF_X1 StateReg_s_current_state_reg_19__FF_FF ( .D(AddRoundKeyOutput[19]), 
        .CK(clk), .Q(ciphertext[19]), .QN() );
  INV_X1 StateReg_s_current_state_reg_18__U1 ( .A(ciphertext[18]), .ZN(
        StateReg_s_current_state_reg_18__QN) );
  DFF_X1 StateReg_s_current_state_reg_18__FF_FF ( .D(AddRoundKeyOutput[18]), 
        .CK(clk), .Q(ciphertext[18]), .QN() );
  INV_X1 StateReg_s_current_state_reg_17__U1 ( .A(ciphertext[17]), .ZN(
        StateReg_s_current_state_reg_17__QN) );
  DFF_X1 StateReg_s_current_state_reg_17__FF_FF ( .D(AddRoundKeyOutput[17]), 
        .CK(clk), .Q(ciphertext[17]), .QN() );
  INV_X1 StateReg_s_current_state_reg_16__U1 ( .A(ciphertext[16]), .ZN(
        StateReg_s_current_state_reg_16__QN) );
  DFF_X1 StateReg_s_current_state_reg_16__FF_FF ( .D(AddRoundKeyOutput[16]), 
        .CK(clk), .Q(ciphertext[16]), .QN() );
  INV_X1 StateReg_s_current_state_reg_15__U1 ( .A(ciphertext[15]), .ZN(
        StateReg_s_current_state_reg_15__QN) );
  DFF_X1 StateReg_s_current_state_reg_15__FF_FF ( .D(AddRoundKeyOutput[15]), 
        .CK(clk), .Q(ciphertext[15]), .QN() );
  INV_X1 StateReg_s_current_state_reg_14__U1 ( .A(ciphertext[14]), .ZN(
        StateReg_s_current_state_reg_14__QN) );
  DFF_X1 StateReg_s_current_state_reg_14__FF_FF ( .D(AddRoundKeyOutput[14]), 
        .CK(clk), .Q(ciphertext[14]), .QN() );
  INV_X1 StateReg_s_current_state_reg_13__U1 ( .A(ciphertext[13]), .ZN(
        StateReg_s_current_state_reg_13__QN) );
  DFF_X1 StateReg_s_current_state_reg_13__FF_FF ( .D(AddRoundKeyOutput[13]), 
        .CK(clk), .Q(ciphertext[13]), .QN() );
  INV_X1 StateReg_s_current_state_reg_12__U1 ( .A(ciphertext[12]), .ZN(
        StateReg_s_current_state_reg_12__QN) );
  DFF_X1 StateReg_s_current_state_reg_12__FF_FF ( .D(AddRoundKeyOutput[12]), 
        .CK(clk), .Q(ciphertext[12]), .QN() );
  INV_X1 StateReg_s_current_state_reg_11__U1 ( .A(ciphertext[11]), .ZN(
        StateReg_s_current_state_reg_11__QN) );
  DFF_X1 StateReg_s_current_state_reg_11__FF_FF ( .D(AddRoundKeyOutput[11]), 
        .CK(clk), .Q(ciphertext[11]), .QN() );
  INV_X1 StateReg_s_current_state_reg_10__U1 ( .A(ciphertext[10]), .ZN(
        StateReg_s_current_state_reg_10__QN) );
  DFF_X1 StateReg_s_current_state_reg_10__FF_FF ( .D(AddRoundKeyOutput[10]), 
        .CK(clk), .Q(ciphertext[10]), .QN() );
  INV_X1 StateReg_s_current_state_reg_9__U1 ( .A(ciphertext[9]), .ZN(
        StateReg_s_current_state_reg_9__QN) );
  DFF_X1 StateReg_s_current_state_reg_9__FF_FF ( .D(AddRoundKeyOutput[9]), 
        .CK(clk), .Q(ciphertext[9]), .QN() );
  INV_X1 StateReg_s_current_state_reg_8__U1 ( .A(ciphertext[8]), .ZN(
        StateReg_s_current_state_reg_8__QN) );
  DFF_X1 StateReg_s_current_state_reg_8__FF_FF ( .D(AddRoundKeyOutput[8]), 
        .CK(clk), .Q(ciphertext[8]), .QN() );
  INV_X1 StateReg_s_current_state_reg_7__U1 ( .A(ciphertext[7]), .ZN(
        StateReg_s_current_state_reg_7__QN) );
  DFF_X1 StateReg_s_current_state_reg_7__FF_FF ( .D(AddRoundKeyOutput[7]), 
        .CK(clk), .Q(ciphertext[7]), .QN() );
  INV_X1 StateReg_s_current_state_reg_6__U1 ( .A(ciphertext[6]), .ZN(
        StateReg_s_current_state_reg_6__QN) );
  DFF_X1 StateReg_s_current_state_reg_6__FF_FF ( .D(AddRoundKeyOutput[6]), 
        .CK(clk), .Q(ciphertext[6]), .QN() );
  INV_X1 StateReg_s_current_state_reg_5__U1 ( .A(ciphertext[5]), .ZN(
        StateReg_s_current_state_reg_5__QN) );
  DFF_X1 StateReg_s_current_state_reg_5__FF_FF ( .D(AddRoundKeyOutput[5]), 
        .CK(clk), .Q(ciphertext[5]), .QN() );
  INV_X1 StateReg_s_current_state_reg_4__U1 ( .A(ciphertext[4]), .ZN(
        StateReg_s_current_state_reg_4__QN) );
  DFF_X1 StateReg_s_current_state_reg_4__FF_FF ( .D(AddRoundKeyOutput[4]), 
        .CK(clk), .Q(ciphertext[4]), .QN() );
  INV_X1 StateReg_s_current_state_reg_3__U1 ( .A(ciphertext[3]), .ZN(
        StateReg_s_current_state_reg_3__QN) );
  DFF_X1 StateReg_s_current_state_reg_3__FF_FF ( .D(AddRoundKeyOutput[3]), 
        .CK(clk), .Q(ciphertext[3]), .QN() );
  INV_X1 StateReg_s_current_state_reg_2__U1 ( .A(ciphertext[2]), .ZN(
        StateReg_s_current_state_reg_2__QN) );
  DFF_X1 StateReg_s_current_state_reg_2__FF_FF ( .D(AddRoundKeyOutput[2]), 
        .CK(clk), .Q(ciphertext[2]), .QN() );
  INV_X1 StateReg_s_current_state_reg_1__U1 ( .A(ciphertext[1]), .ZN(
        StateReg_s_current_state_reg_1__QN) );
  DFF_X1 StateReg_s_current_state_reg_1__FF_FF ( .D(AddRoundKeyOutput[1]), 
        .CK(clk), .Q(ciphertext[1]), .QN() );
  INV_X1 StateReg_s_current_state_reg_0__U1 ( .A(ciphertext[0]), .ZN(
        StateReg_s_current_state_reg_0__QN) );
  DFF_X1 StateReg_s_current_state_reg_0__FF_FF ( .D(AddRoundKeyOutput[0]), 
        .CK(clk), .Q(ciphertext[0]), .QN() );
  NAND2_X1 SubCellInst_SboxInst_0_U19 ( .A1(SubCellInst_SboxInst_0_n15), .A2(
        SubCellInst_SboxInst_0_n14), .ZN(Feedback[3]) );
  OR2_X1 SubCellInst_SboxInst_0_U18 ( .A1(SubCellInst_SboxInst_0_n13), .A2(
        ciphertext[61]), .ZN(SubCellInst_SboxInst_0_n14) );
  NAND2_X1 SubCellInst_SboxInst_0_U17 ( .A1(SubCellInst_SboxInst_0_n15), .A2(
        SubCellInst_SboxInst_0_n12), .ZN(Feedback[2]) );
  NAND2_X1 SubCellInst_SboxInst_0_U16 ( .A1(SubCellInst_SboxInst_0_n11), .A2(
        ciphertext[61]), .ZN(SubCellInst_SboxInst_0_n12) );
  NAND2_X1 SubCellInst_SboxInst_0_U15 ( .A1(SubCellInst_SboxInst_0_n10), .A2(
        SubCellInst_SboxInst_0_n9), .ZN(SubCellInst_SboxInst_0_n11) );
  NAND2_X1 SubCellInst_SboxInst_0_U14 ( .A1(ciphertext[60]), .A2(ciphertext[63]), .ZN(
        SubCellInst_SboxInst_0_n10) );
  NAND2_X1 SubCellInst_SboxInst_0_U13 ( .A1(SubCellInst_SboxInst_0_n8), .A2(
        SubCellInst_SboxInst_0_n7), .ZN(SubCellInst_SboxInst_0_n15) );
  NAND2_X1 SubCellInst_SboxInst_0_U12 ( .A1(SubCellInst_SboxInst_0_n6), .A2(
        SubCellInst_SboxInst_0_n5), .ZN(Feedback[1]) );
  NAND2_X1 SubCellInst_SboxInst_0_U11 ( .A1(ciphertext[60]), .A2(
        SubCellInst_SboxInst_0_n4), .ZN(SubCellInst_SboxInst_0_n5) );
  NAND2_X1 SubCellInst_SboxInst_0_U10 ( .A1(ciphertext[63]), .A2(
        SubCellInst_SboxInst_0_n9), .ZN(SubCellInst_SboxInst_0_n4) );
  NAND2_X1 SubCellInst_SboxInst_0_U9 ( .A1(ciphertext[62]), .A2(
        SubCellInst_SboxInst_0_n8), .ZN(SubCellInst_SboxInst_0_n6) );
  NOR2_X1 SubCellInst_SboxInst_0_U8 ( .A1(SubCellInst_SboxInst_0_n13), .A2(
        SubCellInst_SboxInst_0_n3), .ZN(Feedback[0]) );
  NOR2_X1 SubCellInst_SboxInst_0_U7 ( .A1(ciphertext[61]), .A2(
        SubCellInst_SboxInst_0_n2), .ZN(SubCellInst_SboxInst_0_n3) );
  NOR2_X1 SubCellInst_SboxInst_0_U6 ( .A1(SubCellInst_SboxInst_0_n7), .A2(
        SubCellInst_SboxInst_0_n1), .ZN(SubCellInst_SboxInst_0_n2) );
  NOR2_X1 SubCellInst_SboxInst_0_U5 ( .A1(ciphertext[62]), .A2(ciphertext[63]), .ZN(
        SubCellInst_SboxInst_0_n1) );
  INV_X1 SubCellInst_SboxInst_0_U4 ( .A(ciphertext[60]), .ZN(
        SubCellInst_SboxInst_0_n7) );
  NOR2_X1 SubCellInst_SboxInst_0_U3 ( .A1(SubCellInst_SboxInst_0_n9), .A2(
        SubCellInst_SboxInst_0_n8), .ZN(SubCellInst_SboxInst_0_n13) );
  INV_X1 SubCellInst_SboxInst_0_U2 ( .A(ciphertext[63]), .ZN(
        SubCellInst_SboxInst_0_n8) );
  INV_X1 SubCellInst_SboxInst_0_U1 ( .A(ciphertext[62]), .ZN(
        SubCellInst_SboxInst_0_n9) );
  NAND2_X1 SubCellInst_SboxInst_1_U19 ( .A1(SubCellInst_SboxInst_1_n15), .A2(
        SubCellInst_SboxInst_1_n14), .ZN(Feedback[7]) );
  OR2_X1 SubCellInst_SboxInst_1_U18 ( .A1(SubCellInst_SboxInst_1_n13), .A2(
        ciphertext[49]), .ZN(SubCellInst_SboxInst_1_n14) );
  NAND2_X1 SubCellInst_SboxInst_1_U17 ( .A1(SubCellInst_SboxInst_1_n15), .A2(
        SubCellInst_SboxInst_1_n12), .ZN(Feedback[6]) );
  NAND2_X1 SubCellInst_SboxInst_1_U16 ( .A1(SubCellInst_SboxInst_1_n11), .A2(
        ciphertext[49]), .ZN(SubCellInst_SboxInst_1_n12) );
  NAND2_X1 SubCellInst_SboxInst_1_U15 ( .A1(SubCellInst_SboxInst_1_n10), .A2(
        SubCellInst_SboxInst_1_n9), .ZN(SubCellInst_SboxInst_1_n11) );
  NAND2_X1 SubCellInst_SboxInst_1_U14 ( .A1(ciphertext[48]), .A2(ciphertext[51]), .ZN(
        SubCellInst_SboxInst_1_n10) );
  NAND2_X1 SubCellInst_SboxInst_1_U13 ( .A1(SubCellInst_SboxInst_1_n8), .A2(
        SubCellInst_SboxInst_1_n7), .ZN(SubCellInst_SboxInst_1_n15) );
  NAND2_X1 SubCellInst_SboxInst_1_U12 ( .A1(SubCellInst_SboxInst_1_n6), .A2(
        SubCellInst_SboxInst_1_n5), .ZN(Feedback[5]) );
  NAND2_X1 SubCellInst_SboxInst_1_U11 ( .A1(ciphertext[48]), .A2(
        SubCellInst_SboxInst_1_n4), .ZN(SubCellInst_SboxInst_1_n5) );
  NAND2_X1 SubCellInst_SboxInst_1_U10 ( .A1(ciphertext[51]), .A2(
        SubCellInst_SboxInst_1_n9), .ZN(SubCellInst_SboxInst_1_n4) );
  NAND2_X1 SubCellInst_SboxInst_1_U9 ( .A1(ciphertext[50]), .A2(
        SubCellInst_SboxInst_1_n8), .ZN(SubCellInst_SboxInst_1_n6) );
  NOR2_X1 SubCellInst_SboxInst_1_U8 ( .A1(SubCellInst_SboxInst_1_n13), .A2(
        SubCellInst_SboxInst_1_n3), .ZN(Feedback[4]) );
  NOR2_X1 SubCellInst_SboxInst_1_U7 ( .A1(ciphertext[49]), .A2(
        SubCellInst_SboxInst_1_n2), .ZN(SubCellInst_SboxInst_1_n3) );
  NOR2_X1 SubCellInst_SboxInst_1_U6 ( .A1(SubCellInst_SboxInst_1_n7), .A2(
        SubCellInst_SboxInst_1_n1), .ZN(SubCellInst_SboxInst_1_n2) );
  NOR2_X1 SubCellInst_SboxInst_1_U5 ( .A1(ciphertext[50]), .A2(ciphertext[51]), .ZN(
        SubCellInst_SboxInst_1_n1) );
  INV_X1 SubCellInst_SboxInst_1_U4 ( .A(ciphertext[48]), .ZN(
        SubCellInst_SboxInst_1_n7) );
  NOR2_X1 SubCellInst_SboxInst_1_U3 ( .A1(SubCellInst_SboxInst_1_n9), .A2(
        SubCellInst_SboxInst_1_n8), .ZN(SubCellInst_SboxInst_1_n13) );
  INV_X1 SubCellInst_SboxInst_1_U2 ( .A(ciphertext[51]), .ZN(
        SubCellInst_SboxInst_1_n8) );
  INV_X1 SubCellInst_SboxInst_1_U1 ( .A(ciphertext[50]), .ZN(
        SubCellInst_SboxInst_1_n9) );
  NAND2_X1 SubCellInst_SboxInst_2_U19 ( .A1(SubCellInst_SboxInst_2_n15), .A2(
        SubCellInst_SboxInst_2_n14), .ZN(Feedback[11]) );
  OR2_X1 SubCellInst_SboxInst_2_U18 ( .A1(SubCellInst_SboxInst_2_n13), .A2(
        ciphertext[53]), .ZN(SubCellInst_SboxInst_2_n14) );
  NAND2_X1 SubCellInst_SboxInst_2_U17 ( .A1(SubCellInst_SboxInst_2_n15), .A2(
        SubCellInst_SboxInst_2_n12), .ZN(Feedback[10]) );
  NAND2_X1 SubCellInst_SboxInst_2_U16 ( .A1(SubCellInst_SboxInst_2_n11), .A2(
        ciphertext[53]), .ZN(SubCellInst_SboxInst_2_n12) );
  NAND2_X1 SubCellInst_SboxInst_2_U15 ( .A1(SubCellInst_SboxInst_2_n10), .A2(
        SubCellInst_SboxInst_2_n9), .ZN(SubCellInst_SboxInst_2_n11) );
  NAND2_X1 SubCellInst_SboxInst_2_U14 ( .A1(ciphertext[52]), .A2(ciphertext[55]), .ZN(
        SubCellInst_SboxInst_2_n10) );
  NAND2_X1 SubCellInst_SboxInst_2_U13 ( .A1(SubCellInst_SboxInst_2_n8), .A2(
        SubCellInst_SboxInst_2_n7), .ZN(SubCellInst_SboxInst_2_n15) );
  NAND2_X1 SubCellInst_SboxInst_2_U12 ( .A1(SubCellInst_SboxInst_2_n6), .A2(
        SubCellInst_SboxInst_2_n5), .ZN(Feedback[9]) );
  NAND2_X1 SubCellInst_SboxInst_2_U11 ( .A1(ciphertext[52]), .A2(
        SubCellInst_SboxInst_2_n4), .ZN(SubCellInst_SboxInst_2_n5) );
  NAND2_X1 SubCellInst_SboxInst_2_U10 ( .A1(ciphertext[55]), .A2(
        SubCellInst_SboxInst_2_n9), .ZN(SubCellInst_SboxInst_2_n4) );
  NAND2_X1 SubCellInst_SboxInst_2_U9 ( .A1(ciphertext[54]), .A2(
        SubCellInst_SboxInst_2_n8), .ZN(SubCellInst_SboxInst_2_n6) );
  NOR2_X1 SubCellInst_SboxInst_2_U8 ( .A1(SubCellInst_SboxInst_2_n13), .A2(
        SubCellInst_SboxInst_2_n3), .ZN(Feedback[8]) );
  NOR2_X1 SubCellInst_SboxInst_2_U7 ( .A1(ciphertext[53]), .A2(
        SubCellInst_SboxInst_2_n2), .ZN(SubCellInst_SboxInst_2_n3) );
  NOR2_X1 SubCellInst_SboxInst_2_U6 ( .A1(SubCellInst_SboxInst_2_n7), .A2(
        SubCellInst_SboxInst_2_n1), .ZN(SubCellInst_SboxInst_2_n2) );
  NOR2_X1 SubCellInst_SboxInst_2_U5 ( .A1(ciphertext[54]), .A2(ciphertext[55]), .ZN(
        SubCellInst_SboxInst_2_n1) );
  INV_X1 SubCellInst_SboxInst_2_U4 ( .A(ciphertext[52]), .ZN(
        SubCellInst_SboxInst_2_n7) );
  NOR2_X1 SubCellInst_SboxInst_2_U3 ( .A1(SubCellInst_SboxInst_2_n9), .A2(
        SubCellInst_SboxInst_2_n8), .ZN(SubCellInst_SboxInst_2_n13) );
  INV_X1 SubCellInst_SboxInst_2_U2 ( .A(ciphertext[55]), .ZN(
        SubCellInst_SboxInst_2_n8) );
  INV_X1 SubCellInst_SboxInst_2_U1 ( .A(ciphertext[54]), .ZN(
        SubCellInst_SboxInst_2_n9) );
  NAND2_X1 SubCellInst_SboxInst_3_U19 ( .A1(SubCellInst_SboxInst_3_n15), .A2(
        SubCellInst_SboxInst_3_n14), .ZN(Feedback[15]) );
  OR2_X1 SubCellInst_SboxInst_3_U18 ( .A1(SubCellInst_SboxInst_3_n13), .A2(
        ciphertext[57]), .ZN(SubCellInst_SboxInst_3_n14) );
  NAND2_X1 SubCellInst_SboxInst_3_U17 ( .A1(SubCellInst_SboxInst_3_n15), .A2(
        SubCellInst_SboxInst_3_n12), .ZN(Feedback[14]) );
  NAND2_X1 SubCellInst_SboxInst_3_U16 ( .A1(SubCellInst_SboxInst_3_n11), .A2(
        ciphertext[57]), .ZN(SubCellInst_SboxInst_3_n12) );
  NAND2_X1 SubCellInst_SboxInst_3_U15 ( .A1(SubCellInst_SboxInst_3_n10), .A2(
        SubCellInst_SboxInst_3_n9), .ZN(SubCellInst_SboxInst_3_n11) );
  NAND2_X1 SubCellInst_SboxInst_3_U14 ( .A1(ciphertext[56]), .A2(ciphertext[59]), .ZN(
        SubCellInst_SboxInst_3_n10) );
  NAND2_X1 SubCellInst_SboxInst_3_U13 ( .A1(SubCellInst_SboxInst_3_n8), .A2(
        SubCellInst_SboxInst_3_n7), .ZN(SubCellInst_SboxInst_3_n15) );
  NAND2_X1 SubCellInst_SboxInst_3_U12 ( .A1(SubCellInst_SboxInst_3_n6), .A2(
        SubCellInst_SboxInst_3_n5), .ZN(Feedback[13]) );
  NAND2_X1 SubCellInst_SboxInst_3_U11 ( .A1(ciphertext[56]), .A2(
        SubCellInst_SboxInst_3_n4), .ZN(SubCellInst_SboxInst_3_n5) );
  NAND2_X1 SubCellInst_SboxInst_3_U10 ( .A1(ciphertext[59]), .A2(
        SubCellInst_SboxInst_3_n9), .ZN(SubCellInst_SboxInst_3_n4) );
  NAND2_X1 SubCellInst_SboxInst_3_U9 ( .A1(ciphertext[58]), .A2(
        SubCellInst_SboxInst_3_n8), .ZN(SubCellInst_SboxInst_3_n6) );
  NOR2_X1 SubCellInst_SboxInst_3_U8 ( .A1(SubCellInst_SboxInst_3_n13), .A2(
        SubCellInst_SboxInst_3_n3), .ZN(Feedback[12]) );
  NOR2_X1 SubCellInst_SboxInst_3_U7 ( .A1(ciphertext[57]), .A2(
        SubCellInst_SboxInst_3_n2), .ZN(SubCellInst_SboxInst_3_n3) );
  NOR2_X1 SubCellInst_SboxInst_3_U6 ( .A1(SubCellInst_SboxInst_3_n7), .A2(
        SubCellInst_SboxInst_3_n1), .ZN(SubCellInst_SboxInst_3_n2) );
  NOR2_X1 SubCellInst_SboxInst_3_U5 ( .A1(ciphertext[58]), .A2(ciphertext[59]), .ZN(
        SubCellInst_SboxInst_3_n1) );
  INV_X1 SubCellInst_SboxInst_3_U4 ( .A(ciphertext[56]), .ZN(
        SubCellInst_SboxInst_3_n7) );
  NOR2_X1 SubCellInst_SboxInst_3_U3 ( .A1(SubCellInst_SboxInst_3_n9), .A2(
        SubCellInst_SboxInst_3_n8), .ZN(SubCellInst_SboxInst_3_n13) );
  INV_X1 SubCellInst_SboxInst_3_U2 ( .A(ciphertext[59]), .ZN(
        SubCellInst_SboxInst_3_n8) );
  INV_X1 SubCellInst_SboxInst_3_U1 ( .A(ciphertext[58]), .ZN(
        SubCellInst_SboxInst_3_n9) );
  NAND2_X1 SubCellInst_SboxInst_4_U19 ( .A1(SubCellInst_SboxInst_4_n15), .A2(
        SubCellInst_SboxInst_4_n14), .ZN(Feedback[19]) );
  OR2_X1 SubCellInst_SboxInst_4_U18 ( .A1(SubCellInst_SboxInst_4_n13), .A2(
        ciphertext[33]), .ZN(SubCellInst_SboxInst_4_n14) );
  NAND2_X1 SubCellInst_SboxInst_4_U17 ( .A1(SubCellInst_SboxInst_4_n15), .A2(
        SubCellInst_SboxInst_4_n12), .ZN(Feedback[18]) );
  NAND2_X1 SubCellInst_SboxInst_4_U16 ( .A1(SubCellInst_SboxInst_4_n11), .A2(
        ciphertext[33]), .ZN(SubCellInst_SboxInst_4_n12) );
  NAND2_X1 SubCellInst_SboxInst_4_U15 ( .A1(SubCellInst_SboxInst_4_n10), .A2(
        SubCellInst_SboxInst_4_n9), .ZN(SubCellInst_SboxInst_4_n11) );
  NAND2_X1 SubCellInst_SboxInst_4_U14 ( .A1(ciphertext[32]), .A2(ciphertext[35]), .ZN(
        SubCellInst_SboxInst_4_n10) );
  NAND2_X1 SubCellInst_SboxInst_4_U13 ( .A1(SubCellInst_SboxInst_4_n8), .A2(
        SubCellInst_SboxInst_4_n7), .ZN(SubCellInst_SboxInst_4_n15) );
  NAND2_X1 SubCellInst_SboxInst_4_U12 ( .A1(SubCellInst_SboxInst_4_n6), .A2(
        SubCellInst_SboxInst_4_n5), .ZN(Feedback[17]) );
  NAND2_X1 SubCellInst_SboxInst_4_U11 ( .A1(ciphertext[32]), .A2(
        SubCellInst_SboxInst_4_n4), .ZN(SubCellInst_SboxInst_4_n5) );
  NAND2_X1 SubCellInst_SboxInst_4_U10 ( .A1(ciphertext[35]), .A2(
        SubCellInst_SboxInst_4_n9), .ZN(SubCellInst_SboxInst_4_n4) );
  NAND2_X1 SubCellInst_SboxInst_4_U9 ( .A1(ciphertext[34]), .A2(
        SubCellInst_SboxInst_4_n8), .ZN(SubCellInst_SboxInst_4_n6) );
  NOR2_X1 SubCellInst_SboxInst_4_U8 ( .A1(SubCellInst_SboxInst_4_n13), .A2(
        SubCellInst_SboxInst_4_n3), .ZN(Feedback[16]) );
  NOR2_X1 SubCellInst_SboxInst_4_U7 ( .A1(ciphertext[33]), .A2(
        SubCellInst_SboxInst_4_n2), .ZN(SubCellInst_SboxInst_4_n3) );
  NOR2_X1 SubCellInst_SboxInst_4_U6 ( .A1(SubCellInst_SboxInst_4_n7), .A2(
        SubCellInst_SboxInst_4_n1), .ZN(SubCellInst_SboxInst_4_n2) );
  NOR2_X1 SubCellInst_SboxInst_4_U5 ( .A1(ciphertext[34]), .A2(ciphertext[35]), .ZN(
        SubCellInst_SboxInst_4_n1) );
  INV_X1 SubCellInst_SboxInst_4_U4 ( .A(ciphertext[32]), .ZN(
        SubCellInst_SboxInst_4_n7) );
  NOR2_X1 SubCellInst_SboxInst_4_U3 ( .A1(SubCellInst_SboxInst_4_n9), .A2(
        SubCellInst_SboxInst_4_n8), .ZN(SubCellInst_SboxInst_4_n13) );
  INV_X1 SubCellInst_SboxInst_4_U2 ( .A(ciphertext[35]), .ZN(
        SubCellInst_SboxInst_4_n8) );
  INV_X1 SubCellInst_SboxInst_4_U1 ( .A(ciphertext[34]), .ZN(
        SubCellInst_SboxInst_4_n9) );
  NAND2_X1 SubCellInst_SboxInst_5_U19 ( .A1(SubCellInst_SboxInst_5_n15), .A2(
        SubCellInst_SboxInst_5_n14), .ZN(Feedback[23]) );
  OR2_X1 SubCellInst_SboxInst_5_U18 ( .A1(SubCellInst_SboxInst_5_n13), .A2(
        ciphertext[45]), .ZN(SubCellInst_SboxInst_5_n14) );
  NAND2_X1 SubCellInst_SboxInst_5_U17 ( .A1(SubCellInst_SboxInst_5_n15), .A2(
        SubCellInst_SboxInst_5_n12), .ZN(Feedback[22]) );
  NAND2_X1 SubCellInst_SboxInst_5_U16 ( .A1(SubCellInst_SboxInst_5_n11), .A2(
        ciphertext[45]), .ZN(SubCellInst_SboxInst_5_n12) );
  NAND2_X1 SubCellInst_SboxInst_5_U15 ( .A1(SubCellInst_SboxInst_5_n10), .A2(
        SubCellInst_SboxInst_5_n9), .ZN(SubCellInst_SboxInst_5_n11) );
  NAND2_X1 SubCellInst_SboxInst_5_U14 ( .A1(ciphertext[44]), .A2(ciphertext[47]), .ZN(
        SubCellInst_SboxInst_5_n10) );
  NAND2_X1 SubCellInst_SboxInst_5_U13 ( .A1(SubCellInst_SboxInst_5_n8), .A2(
        SubCellInst_SboxInst_5_n7), .ZN(SubCellInst_SboxInst_5_n15) );
  NAND2_X1 SubCellInst_SboxInst_5_U12 ( .A1(SubCellInst_SboxInst_5_n6), .A2(
        SubCellInst_SboxInst_5_n5), .ZN(Feedback[21]) );
  NAND2_X1 SubCellInst_SboxInst_5_U11 ( .A1(ciphertext[44]), .A2(
        SubCellInst_SboxInst_5_n4), .ZN(SubCellInst_SboxInst_5_n5) );
  NAND2_X1 SubCellInst_SboxInst_5_U10 ( .A1(ciphertext[47]), .A2(
        SubCellInst_SboxInst_5_n9), .ZN(SubCellInst_SboxInst_5_n4) );
  NAND2_X1 SubCellInst_SboxInst_5_U9 ( .A1(ciphertext[46]), .A2(
        SubCellInst_SboxInst_5_n8), .ZN(SubCellInst_SboxInst_5_n6) );
  NOR2_X1 SubCellInst_SboxInst_5_U8 ( .A1(SubCellInst_SboxInst_5_n13), .A2(
        SubCellInst_SboxInst_5_n3), .ZN(Feedback[20]) );
  NOR2_X1 SubCellInst_SboxInst_5_U7 ( .A1(ciphertext[45]), .A2(
        SubCellInst_SboxInst_5_n2), .ZN(SubCellInst_SboxInst_5_n3) );
  NOR2_X1 SubCellInst_SboxInst_5_U6 ( .A1(SubCellInst_SboxInst_5_n7), .A2(
        SubCellInst_SboxInst_5_n1), .ZN(SubCellInst_SboxInst_5_n2) );
  NOR2_X1 SubCellInst_SboxInst_5_U5 ( .A1(ciphertext[46]), .A2(ciphertext[47]), .ZN(
        SubCellInst_SboxInst_5_n1) );
  INV_X1 SubCellInst_SboxInst_5_U4 ( .A(ciphertext[44]), .ZN(
        SubCellInst_SboxInst_5_n7) );
  NOR2_X1 SubCellInst_SboxInst_5_U3 ( .A1(SubCellInst_SboxInst_5_n9), .A2(
        SubCellInst_SboxInst_5_n8), .ZN(SubCellInst_SboxInst_5_n13) );
  INV_X1 SubCellInst_SboxInst_5_U2 ( .A(ciphertext[47]), .ZN(
        SubCellInst_SboxInst_5_n8) );
  INV_X1 SubCellInst_SboxInst_5_U1 ( .A(ciphertext[46]), .ZN(
        SubCellInst_SboxInst_5_n9) );
  NAND2_X1 SubCellInst_SboxInst_6_U19 ( .A1(SubCellInst_SboxInst_6_n15), .A2(
        SubCellInst_SboxInst_6_n14), .ZN(Feedback[27]) );
  OR2_X1 SubCellInst_SboxInst_6_U18 ( .A1(SubCellInst_SboxInst_6_n13), .A2(
        ciphertext[41]), .ZN(SubCellInst_SboxInst_6_n14) );
  NAND2_X1 SubCellInst_SboxInst_6_U17 ( .A1(SubCellInst_SboxInst_6_n15), .A2(
        SubCellInst_SboxInst_6_n12), .ZN(Feedback[26]) );
  NAND2_X1 SubCellInst_SboxInst_6_U16 ( .A1(SubCellInst_SboxInst_6_n11), .A2(
        ciphertext[41]), .ZN(SubCellInst_SboxInst_6_n12) );
  NAND2_X1 SubCellInst_SboxInst_6_U15 ( .A1(SubCellInst_SboxInst_6_n10), .A2(
        SubCellInst_SboxInst_6_n9), .ZN(SubCellInst_SboxInst_6_n11) );
  NAND2_X1 SubCellInst_SboxInst_6_U14 ( .A1(ciphertext[40]), .A2(ciphertext[43]), .ZN(
        SubCellInst_SboxInst_6_n10) );
  NAND2_X1 SubCellInst_SboxInst_6_U13 ( .A1(SubCellInst_SboxInst_6_n8), .A2(
        SubCellInst_SboxInst_6_n7), .ZN(SubCellInst_SboxInst_6_n15) );
  NAND2_X1 SubCellInst_SboxInst_6_U12 ( .A1(SubCellInst_SboxInst_6_n6), .A2(
        SubCellInst_SboxInst_6_n5), .ZN(Feedback[25]) );
  NAND2_X1 SubCellInst_SboxInst_6_U11 ( .A1(ciphertext[40]), .A2(
        SubCellInst_SboxInst_6_n4), .ZN(SubCellInst_SboxInst_6_n5) );
  NAND2_X1 SubCellInst_SboxInst_6_U10 ( .A1(ciphertext[43]), .A2(
        SubCellInst_SboxInst_6_n9), .ZN(SubCellInst_SboxInst_6_n4) );
  NAND2_X1 SubCellInst_SboxInst_6_U9 ( .A1(ciphertext[42]), .A2(
        SubCellInst_SboxInst_6_n8), .ZN(SubCellInst_SboxInst_6_n6) );
  NOR2_X1 SubCellInst_SboxInst_6_U8 ( .A1(SubCellInst_SboxInst_6_n13), .A2(
        SubCellInst_SboxInst_6_n3), .ZN(Feedback[24]) );
  NOR2_X1 SubCellInst_SboxInst_6_U7 ( .A1(ciphertext[41]), .A2(
        SubCellInst_SboxInst_6_n2), .ZN(SubCellInst_SboxInst_6_n3) );
  NOR2_X1 SubCellInst_SboxInst_6_U6 ( .A1(SubCellInst_SboxInst_6_n7), .A2(
        SubCellInst_SboxInst_6_n1), .ZN(SubCellInst_SboxInst_6_n2) );
  NOR2_X1 SubCellInst_SboxInst_6_U5 ( .A1(ciphertext[42]), .A2(ciphertext[43]), .ZN(
        SubCellInst_SboxInst_6_n1) );
  INV_X1 SubCellInst_SboxInst_6_U4 ( .A(ciphertext[40]), .ZN(
        SubCellInst_SboxInst_6_n7) );
  NOR2_X1 SubCellInst_SboxInst_6_U3 ( .A1(SubCellInst_SboxInst_6_n9), .A2(
        SubCellInst_SboxInst_6_n8), .ZN(SubCellInst_SboxInst_6_n13) );
  INV_X1 SubCellInst_SboxInst_6_U2 ( .A(ciphertext[43]), .ZN(
        SubCellInst_SboxInst_6_n8) );
  INV_X1 SubCellInst_SboxInst_6_U1 ( .A(ciphertext[42]), .ZN(
        SubCellInst_SboxInst_6_n9) );
  NAND2_X1 SubCellInst_SboxInst_7_U19 ( .A1(SubCellInst_SboxInst_7_n15), .A2(
        SubCellInst_SboxInst_7_n14), .ZN(Feedback[31]) );
  OR2_X1 SubCellInst_SboxInst_7_U18 ( .A1(SubCellInst_SboxInst_7_n13), .A2(
        ciphertext[37]), .ZN(SubCellInst_SboxInst_7_n14) );
  NAND2_X1 SubCellInst_SboxInst_7_U17 ( .A1(SubCellInst_SboxInst_7_n15), .A2(
        SubCellInst_SboxInst_7_n12), .ZN(Feedback[30]) );
  NAND2_X1 SubCellInst_SboxInst_7_U16 ( .A1(SubCellInst_SboxInst_7_n11), .A2(
        ciphertext[37]), .ZN(SubCellInst_SboxInst_7_n12) );
  NAND2_X1 SubCellInst_SboxInst_7_U15 ( .A1(SubCellInst_SboxInst_7_n10), .A2(
        SubCellInst_SboxInst_7_n9), .ZN(SubCellInst_SboxInst_7_n11) );
  NAND2_X1 SubCellInst_SboxInst_7_U14 ( .A1(ciphertext[36]), .A2(ciphertext[39]), .ZN(
        SubCellInst_SboxInst_7_n10) );
  NAND2_X1 SubCellInst_SboxInst_7_U13 ( .A1(SubCellInst_SboxInst_7_n8), .A2(
        SubCellInst_SboxInst_7_n7), .ZN(SubCellInst_SboxInst_7_n15) );
  NAND2_X1 SubCellInst_SboxInst_7_U12 ( .A1(SubCellInst_SboxInst_7_n6), .A2(
        SubCellInst_SboxInst_7_n5), .ZN(Feedback[29]) );
  NAND2_X1 SubCellInst_SboxInst_7_U11 ( .A1(ciphertext[36]), .A2(
        SubCellInst_SboxInst_7_n4), .ZN(SubCellInst_SboxInst_7_n5) );
  NAND2_X1 SubCellInst_SboxInst_7_U10 ( .A1(ciphertext[39]), .A2(
        SubCellInst_SboxInst_7_n9), .ZN(SubCellInst_SboxInst_7_n4) );
  NAND2_X1 SubCellInst_SboxInst_7_U9 ( .A1(ciphertext[38]), .A2(
        SubCellInst_SboxInst_7_n8), .ZN(SubCellInst_SboxInst_7_n6) );
  NOR2_X1 SubCellInst_SboxInst_7_U8 ( .A1(SubCellInst_SboxInst_7_n13), .A2(
        SubCellInst_SboxInst_7_n3), .ZN(Feedback[28]) );
  NOR2_X1 SubCellInst_SboxInst_7_U7 ( .A1(ciphertext[37]), .A2(
        SubCellInst_SboxInst_7_n2), .ZN(SubCellInst_SboxInst_7_n3) );
  NOR2_X1 SubCellInst_SboxInst_7_U6 ( .A1(SubCellInst_SboxInst_7_n7), .A2(
        SubCellInst_SboxInst_7_n1), .ZN(SubCellInst_SboxInst_7_n2) );
  NOR2_X1 SubCellInst_SboxInst_7_U5 ( .A1(ciphertext[38]), .A2(ciphertext[39]), .ZN(
        SubCellInst_SboxInst_7_n1) );
  INV_X1 SubCellInst_SboxInst_7_U4 ( .A(ciphertext[36]), .ZN(
        SubCellInst_SboxInst_7_n7) );
  NOR2_X1 SubCellInst_SboxInst_7_U3 ( .A1(SubCellInst_SboxInst_7_n9), .A2(
        SubCellInst_SboxInst_7_n8), .ZN(SubCellInst_SboxInst_7_n13) );
  INV_X1 SubCellInst_SboxInst_7_U2 ( .A(ciphertext[39]), .ZN(
        SubCellInst_SboxInst_7_n8) );
  INV_X1 SubCellInst_SboxInst_7_U1 ( .A(ciphertext[38]), .ZN(
        SubCellInst_SboxInst_7_n9) );
  NAND2_X1 SubCellInst_SboxInst_8_U19 ( .A1(SubCellInst_SboxInst_8_n15), .A2(
        SubCellInst_SboxInst_8_n14), .ZN(Feedback[35]) );
  OR2_X1 SubCellInst_SboxInst_8_U18 ( .A1(SubCellInst_SboxInst_8_n13), .A2(
        ciphertext[17]), .ZN(SubCellInst_SboxInst_8_n14) );
  NAND2_X1 SubCellInst_SboxInst_8_U17 ( .A1(SubCellInst_SboxInst_8_n15), .A2(
        SubCellInst_SboxInst_8_n12), .ZN(Feedback[34]) );
  NAND2_X1 SubCellInst_SboxInst_8_U16 ( .A1(SubCellInst_SboxInst_8_n11), .A2(
        ciphertext[17]), .ZN(SubCellInst_SboxInst_8_n12) );
  NAND2_X1 SubCellInst_SboxInst_8_U15 ( .A1(SubCellInst_SboxInst_8_n10), .A2(
        SubCellInst_SboxInst_8_n9), .ZN(SubCellInst_SboxInst_8_n11) );
  NAND2_X1 SubCellInst_SboxInst_8_U14 ( .A1(ciphertext[16]), .A2(ciphertext[19]), .ZN(
        SubCellInst_SboxInst_8_n10) );
  NAND2_X1 SubCellInst_SboxInst_8_U13 ( .A1(SubCellInst_SboxInst_8_n8), .A2(
        SubCellInst_SboxInst_8_n7), .ZN(SubCellInst_SboxInst_8_n15) );
  NAND2_X1 SubCellInst_SboxInst_8_U12 ( .A1(SubCellInst_SboxInst_8_n6), .A2(
        SubCellInst_SboxInst_8_n5), .ZN(Feedback[33]) );
  NAND2_X1 SubCellInst_SboxInst_8_U11 ( .A1(ciphertext[16]), .A2(
        SubCellInst_SboxInst_8_n4), .ZN(SubCellInst_SboxInst_8_n5) );
  NAND2_X1 SubCellInst_SboxInst_8_U10 ( .A1(ciphertext[19]), .A2(
        SubCellInst_SboxInst_8_n9), .ZN(SubCellInst_SboxInst_8_n4) );
  NAND2_X1 SubCellInst_SboxInst_8_U9 ( .A1(ciphertext[18]), .A2(
        SubCellInst_SboxInst_8_n8), .ZN(SubCellInst_SboxInst_8_n6) );
  NOR2_X1 SubCellInst_SboxInst_8_U8 ( .A1(SubCellInst_SboxInst_8_n13), .A2(
        SubCellInst_SboxInst_8_n3), .ZN(Feedback[32]) );
  NOR2_X1 SubCellInst_SboxInst_8_U7 ( .A1(ciphertext[17]), .A2(
        SubCellInst_SboxInst_8_n2), .ZN(SubCellInst_SboxInst_8_n3) );
  NOR2_X1 SubCellInst_SboxInst_8_U6 ( .A1(SubCellInst_SboxInst_8_n7), .A2(
        SubCellInst_SboxInst_8_n1), .ZN(SubCellInst_SboxInst_8_n2) );
  NOR2_X1 SubCellInst_SboxInst_8_U5 ( .A1(ciphertext[18]), .A2(ciphertext[19]), .ZN(
        SubCellInst_SboxInst_8_n1) );
  INV_X1 SubCellInst_SboxInst_8_U4 ( .A(ciphertext[16]), .ZN(
        SubCellInst_SboxInst_8_n7) );
  NOR2_X1 SubCellInst_SboxInst_8_U3 ( .A1(SubCellInst_SboxInst_8_n9), .A2(
        SubCellInst_SboxInst_8_n8), .ZN(SubCellInst_SboxInst_8_n13) );
  INV_X1 SubCellInst_SboxInst_8_U2 ( .A(ciphertext[19]), .ZN(
        SubCellInst_SboxInst_8_n8) );
  INV_X1 SubCellInst_SboxInst_8_U1 ( .A(ciphertext[18]), .ZN(
        SubCellInst_SboxInst_8_n9) );
  NAND2_X1 SubCellInst_SboxInst_9_U19 ( .A1(SubCellInst_SboxInst_9_n15), .A2(
        SubCellInst_SboxInst_9_n14), .ZN(Feedback[39]) );
  OR2_X1 SubCellInst_SboxInst_9_U18 ( .A1(SubCellInst_SboxInst_9_n13), .A2(
        ciphertext[29]), .ZN(SubCellInst_SboxInst_9_n14) );
  NAND2_X1 SubCellInst_SboxInst_9_U17 ( .A1(SubCellInst_SboxInst_9_n15), .A2(
        SubCellInst_SboxInst_9_n12), .ZN(Feedback[38]) );
  NAND2_X1 SubCellInst_SboxInst_9_U16 ( .A1(SubCellInst_SboxInst_9_n11), .A2(
        ciphertext[29]), .ZN(SubCellInst_SboxInst_9_n12) );
  NAND2_X1 SubCellInst_SboxInst_9_U15 ( .A1(SubCellInst_SboxInst_9_n10), .A2(
        SubCellInst_SboxInst_9_n9), .ZN(SubCellInst_SboxInst_9_n11) );
  NAND2_X1 SubCellInst_SboxInst_9_U14 ( .A1(ciphertext[28]), .A2(ciphertext[31]), .ZN(
        SubCellInst_SboxInst_9_n10) );
  NAND2_X1 SubCellInst_SboxInst_9_U13 ( .A1(SubCellInst_SboxInst_9_n8), .A2(
        SubCellInst_SboxInst_9_n7), .ZN(SubCellInst_SboxInst_9_n15) );
  NAND2_X1 SubCellInst_SboxInst_9_U12 ( .A1(SubCellInst_SboxInst_9_n6), .A2(
        SubCellInst_SboxInst_9_n5), .ZN(Feedback[37]) );
  NAND2_X1 SubCellInst_SboxInst_9_U11 ( .A1(ciphertext[28]), .A2(
        SubCellInst_SboxInst_9_n4), .ZN(SubCellInst_SboxInst_9_n5) );
  NAND2_X1 SubCellInst_SboxInst_9_U10 ( .A1(ciphertext[31]), .A2(
        SubCellInst_SboxInst_9_n9), .ZN(SubCellInst_SboxInst_9_n4) );
  NAND2_X1 SubCellInst_SboxInst_9_U9 ( .A1(ciphertext[30]), .A2(
        SubCellInst_SboxInst_9_n8), .ZN(SubCellInst_SboxInst_9_n6) );
  NOR2_X1 SubCellInst_SboxInst_9_U8 ( .A1(SubCellInst_SboxInst_9_n13), .A2(
        SubCellInst_SboxInst_9_n3), .ZN(Feedback[36]) );
  NOR2_X1 SubCellInst_SboxInst_9_U7 ( .A1(ciphertext[29]), .A2(
        SubCellInst_SboxInst_9_n2), .ZN(SubCellInst_SboxInst_9_n3) );
  NOR2_X1 SubCellInst_SboxInst_9_U6 ( .A1(SubCellInst_SboxInst_9_n7), .A2(
        SubCellInst_SboxInst_9_n1), .ZN(SubCellInst_SboxInst_9_n2) );
  NOR2_X1 SubCellInst_SboxInst_9_U5 ( .A1(ciphertext[30]), .A2(ciphertext[31]), .ZN(
        SubCellInst_SboxInst_9_n1) );
  INV_X1 SubCellInst_SboxInst_9_U4 ( .A(ciphertext[28]), .ZN(
        SubCellInst_SboxInst_9_n7) );
  NOR2_X1 SubCellInst_SboxInst_9_U3 ( .A1(SubCellInst_SboxInst_9_n9), .A2(
        SubCellInst_SboxInst_9_n8), .ZN(SubCellInst_SboxInst_9_n13) );
  INV_X1 SubCellInst_SboxInst_9_U2 ( .A(ciphertext[31]), .ZN(
        SubCellInst_SboxInst_9_n8) );
  INV_X1 SubCellInst_SboxInst_9_U1 ( .A(ciphertext[30]), .ZN(
        SubCellInst_SboxInst_9_n9) );
  NAND2_X1 SubCellInst_SboxInst_10_U19 ( .A1(SubCellInst_SboxInst_10_n15), 
        .A2(SubCellInst_SboxInst_10_n14), .ZN(Feedback[43]) );
  OR2_X1 SubCellInst_SboxInst_10_U18 ( .A1(SubCellInst_SboxInst_10_n13), .A2(
        ciphertext[25]), .ZN(SubCellInst_SboxInst_10_n14) );
  NAND2_X1 SubCellInst_SboxInst_10_U17 ( .A1(SubCellInst_SboxInst_10_n15), 
        .A2(SubCellInst_SboxInst_10_n12), .ZN(Feedback[42]) );
  NAND2_X1 SubCellInst_SboxInst_10_U16 ( .A1(SubCellInst_SboxInst_10_n11), 
        .A2(ciphertext[25]), .ZN(SubCellInst_SboxInst_10_n12) );
  NAND2_X1 SubCellInst_SboxInst_10_U15 ( .A1(SubCellInst_SboxInst_10_n10), 
        .A2(SubCellInst_SboxInst_10_n9), .ZN(SubCellInst_SboxInst_10_n11) );
  NAND2_X1 SubCellInst_SboxInst_10_U14 ( .A1(ciphertext[24]), .A2(ciphertext[27]), 
        .ZN(SubCellInst_SboxInst_10_n10) );
  NAND2_X1 SubCellInst_SboxInst_10_U13 ( .A1(SubCellInst_SboxInst_10_n8), .A2(
        SubCellInst_SboxInst_10_n7), .ZN(SubCellInst_SboxInst_10_n15) );
  NAND2_X1 SubCellInst_SboxInst_10_U12 ( .A1(SubCellInst_SboxInst_10_n6), .A2(
        SubCellInst_SboxInst_10_n5), .ZN(Feedback[41]) );
  NAND2_X1 SubCellInst_SboxInst_10_U11 ( .A1(ciphertext[24]), .A2(
        SubCellInst_SboxInst_10_n4), .ZN(SubCellInst_SboxInst_10_n5) );
  NAND2_X1 SubCellInst_SboxInst_10_U10 ( .A1(ciphertext[27]), .A2(
        SubCellInst_SboxInst_10_n9), .ZN(SubCellInst_SboxInst_10_n4) );
  NAND2_X1 SubCellInst_SboxInst_10_U9 ( .A1(ciphertext[26]), .A2(
        SubCellInst_SboxInst_10_n8), .ZN(SubCellInst_SboxInst_10_n6) );
  NOR2_X1 SubCellInst_SboxInst_10_U8 ( .A1(SubCellInst_SboxInst_10_n13), .A2(
        SubCellInst_SboxInst_10_n3), .ZN(Feedback[40]) );
  NOR2_X1 SubCellInst_SboxInst_10_U7 ( .A1(ciphertext[25]), .A2(
        SubCellInst_SboxInst_10_n2), .ZN(SubCellInst_SboxInst_10_n3) );
  NOR2_X1 SubCellInst_SboxInst_10_U6 ( .A1(SubCellInst_SboxInst_10_n7), .A2(
        SubCellInst_SboxInst_10_n1), .ZN(SubCellInst_SboxInst_10_n2) );
  NOR2_X1 SubCellInst_SboxInst_10_U5 ( .A1(ciphertext[26]), .A2(ciphertext[27]), .ZN(
        SubCellInst_SboxInst_10_n1) );
  INV_X1 SubCellInst_SboxInst_10_U4 ( .A(ciphertext[24]), .ZN(
        SubCellInst_SboxInst_10_n7) );
  NOR2_X1 SubCellInst_SboxInst_10_U3 ( .A1(SubCellInst_SboxInst_10_n9), .A2(
        SubCellInst_SboxInst_10_n8), .ZN(SubCellInst_SboxInst_10_n13) );
  INV_X1 SubCellInst_SboxInst_10_U2 ( .A(ciphertext[27]), .ZN(
        SubCellInst_SboxInst_10_n8) );
  INV_X1 SubCellInst_SboxInst_10_U1 ( .A(ciphertext[26]), .ZN(
        SubCellInst_SboxInst_10_n9) );
  NAND2_X1 SubCellInst_SboxInst_11_U19 ( .A1(SubCellInst_SboxInst_11_n15), 
        .A2(SubCellInst_SboxInst_11_n14), .ZN(Feedback[47]) );
  OR2_X1 SubCellInst_SboxInst_11_U18 ( .A1(SubCellInst_SboxInst_11_n13), .A2(
        ciphertext[21]), .ZN(SubCellInst_SboxInst_11_n14) );
  NAND2_X1 SubCellInst_SboxInst_11_U17 ( .A1(SubCellInst_SboxInst_11_n15), 
        .A2(SubCellInst_SboxInst_11_n12), .ZN(Feedback[46]) );
  NAND2_X1 SubCellInst_SboxInst_11_U16 ( .A1(SubCellInst_SboxInst_11_n11), 
        .A2(ciphertext[21]), .ZN(SubCellInst_SboxInst_11_n12) );
  NAND2_X1 SubCellInst_SboxInst_11_U15 ( .A1(SubCellInst_SboxInst_11_n10), 
        .A2(SubCellInst_SboxInst_11_n9), .ZN(SubCellInst_SboxInst_11_n11) );
  NAND2_X1 SubCellInst_SboxInst_11_U14 ( .A1(ciphertext[20]), .A2(ciphertext[23]), 
        .ZN(SubCellInst_SboxInst_11_n10) );
  NAND2_X1 SubCellInst_SboxInst_11_U13 ( .A1(SubCellInst_SboxInst_11_n8), .A2(
        SubCellInst_SboxInst_11_n7), .ZN(SubCellInst_SboxInst_11_n15) );
  NAND2_X1 SubCellInst_SboxInst_11_U12 ( .A1(SubCellInst_SboxInst_11_n6), .A2(
        SubCellInst_SboxInst_11_n5), .ZN(Feedback[45]) );
  NAND2_X1 SubCellInst_SboxInst_11_U11 ( .A1(ciphertext[20]), .A2(
        SubCellInst_SboxInst_11_n4), .ZN(SubCellInst_SboxInst_11_n5) );
  NAND2_X1 SubCellInst_SboxInst_11_U10 ( .A1(ciphertext[23]), .A2(
        SubCellInst_SboxInst_11_n9), .ZN(SubCellInst_SboxInst_11_n4) );
  NAND2_X1 SubCellInst_SboxInst_11_U9 ( .A1(ciphertext[22]), .A2(
        SubCellInst_SboxInst_11_n8), .ZN(SubCellInst_SboxInst_11_n6) );
  NOR2_X1 SubCellInst_SboxInst_11_U8 ( .A1(SubCellInst_SboxInst_11_n13), .A2(
        SubCellInst_SboxInst_11_n3), .ZN(Feedback[44]) );
  NOR2_X1 SubCellInst_SboxInst_11_U7 ( .A1(ciphertext[21]), .A2(
        SubCellInst_SboxInst_11_n2), .ZN(SubCellInst_SboxInst_11_n3) );
  NOR2_X1 SubCellInst_SboxInst_11_U6 ( .A1(SubCellInst_SboxInst_11_n7), .A2(
        SubCellInst_SboxInst_11_n1), .ZN(SubCellInst_SboxInst_11_n2) );
  NOR2_X1 SubCellInst_SboxInst_11_U5 ( .A1(ciphertext[22]), .A2(ciphertext[23]), .ZN(
        SubCellInst_SboxInst_11_n1) );
  INV_X1 SubCellInst_SboxInst_11_U4 ( .A(ciphertext[20]), .ZN(
        SubCellInst_SboxInst_11_n7) );
  NOR2_X1 SubCellInst_SboxInst_11_U3 ( .A1(SubCellInst_SboxInst_11_n9), .A2(
        SubCellInst_SboxInst_11_n8), .ZN(SubCellInst_SboxInst_11_n13) );
  INV_X1 SubCellInst_SboxInst_11_U2 ( .A(ciphertext[23]), .ZN(
        SubCellInst_SboxInst_11_n8) );
  INV_X1 SubCellInst_SboxInst_11_U1 ( .A(ciphertext[22]), .ZN(
        SubCellInst_SboxInst_11_n9) );
  NAND2_X1 SubCellInst_SboxInst_12_U19 ( .A1(SubCellInst_SboxInst_12_n15), 
        .A2(SubCellInst_SboxInst_12_n14), .ZN(Feedback[51]) );
  OR2_X1 SubCellInst_SboxInst_12_U18 ( .A1(SubCellInst_SboxInst_12_n13), .A2(
        ciphertext[5]), .ZN(SubCellInst_SboxInst_12_n14) );
  NAND2_X1 SubCellInst_SboxInst_12_U17 ( .A1(SubCellInst_SboxInst_12_n15), 
        .A2(SubCellInst_SboxInst_12_n12), .ZN(Feedback[50]) );
  NAND2_X1 SubCellInst_SboxInst_12_U16 ( .A1(SubCellInst_SboxInst_12_n11), 
        .A2(ciphertext[5]), .ZN(SubCellInst_SboxInst_12_n12) );
  NAND2_X1 SubCellInst_SboxInst_12_U15 ( .A1(SubCellInst_SboxInst_12_n10), 
        .A2(SubCellInst_SboxInst_12_n9), .ZN(SubCellInst_SboxInst_12_n11) );
  NAND2_X1 SubCellInst_SboxInst_12_U14 ( .A1(ciphertext[4]), .A2(ciphertext[7]), .ZN(
        SubCellInst_SboxInst_12_n10) );
  NAND2_X1 SubCellInst_SboxInst_12_U13 ( .A1(SubCellInst_SboxInst_12_n8), .A2(
        SubCellInst_SboxInst_12_n7), .ZN(SubCellInst_SboxInst_12_n15) );
  NAND2_X1 SubCellInst_SboxInst_12_U12 ( .A1(SubCellInst_SboxInst_12_n6), .A2(
        SubCellInst_SboxInst_12_n5), .ZN(Feedback[49]) );
  NAND2_X1 SubCellInst_SboxInst_12_U11 ( .A1(ciphertext[4]), .A2(
        SubCellInst_SboxInst_12_n4), .ZN(SubCellInst_SboxInst_12_n5) );
  NAND2_X1 SubCellInst_SboxInst_12_U10 ( .A1(ciphertext[7]), .A2(
        SubCellInst_SboxInst_12_n9), .ZN(SubCellInst_SboxInst_12_n4) );
  NAND2_X1 SubCellInst_SboxInst_12_U9 ( .A1(ciphertext[6]), .A2(
        SubCellInst_SboxInst_12_n8), .ZN(SubCellInst_SboxInst_12_n6) );
  NOR2_X1 SubCellInst_SboxInst_12_U8 ( .A1(SubCellInst_SboxInst_12_n13), .A2(
        SubCellInst_SboxInst_12_n3), .ZN(Feedback[48]) );
  NOR2_X1 SubCellInst_SboxInst_12_U7 ( .A1(ciphertext[5]), .A2(
        SubCellInst_SboxInst_12_n2), .ZN(SubCellInst_SboxInst_12_n3) );
  NOR2_X1 SubCellInst_SboxInst_12_U6 ( .A1(SubCellInst_SboxInst_12_n7), .A2(
        SubCellInst_SboxInst_12_n1), .ZN(SubCellInst_SboxInst_12_n2) );
  NOR2_X1 SubCellInst_SboxInst_12_U5 ( .A1(ciphertext[6]), .A2(ciphertext[7]), .ZN(
        SubCellInst_SboxInst_12_n1) );
  INV_X1 SubCellInst_SboxInst_12_U4 ( .A(ciphertext[4]), .ZN(
        SubCellInst_SboxInst_12_n7) );
  NOR2_X1 SubCellInst_SboxInst_12_U3 ( .A1(SubCellInst_SboxInst_12_n9), .A2(
        SubCellInst_SboxInst_12_n8), .ZN(SubCellInst_SboxInst_12_n13) );
  INV_X1 SubCellInst_SboxInst_12_U2 ( .A(ciphertext[7]), .ZN(
        SubCellInst_SboxInst_12_n8) );
  INV_X1 SubCellInst_SboxInst_12_U1 ( .A(ciphertext[6]), .ZN(
        SubCellInst_SboxInst_12_n9) );
  NAND2_X1 SubCellInst_SboxInst_13_U19 ( .A1(SubCellInst_SboxInst_13_n15), 
        .A2(SubCellInst_SboxInst_13_n14), .ZN(Feedback[55]) );
  OR2_X1 SubCellInst_SboxInst_13_U18 ( .A1(SubCellInst_SboxInst_13_n13), .A2(
        ciphertext[9]), .ZN(SubCellInst_SboxInst_13_n14) );
  NAND2_X1 SubCellInst_SboxInst_13_U17 ( .A1(SubCellInst_SboxInst_13_n15), 
        .A2(SubCellInst_SboxInst_13_n12), .ZN(Feedback[54]) );
  NAND2_X1 SubCellInst_SboxInst_13_U16 ( .A1(SubCellInst_SboxInst_13_n11), 
        .A2(ciphertext[9]), .ZN(SubCellInst_SboxInst_13_n12) );
  NAND2_X1 SubCellInst_SboxInst_13_U15 ( .A1(SubCellInst_SboxInst_13_n10), 
        .A2(SubCellInst_SboxInst_13_n9), .ZN(SubCellInst_SboxInst_13_n11) );
  NAND2_X1 SubCellInst_SboxInst_13_U14 ( .A1(ciphertext[8]), .A2(ciphertext[11]), .ZN(
        SubCellInst_SboxInst_13_n10) );
  NAND2_X1 SubCellInst_SboxInst_13_U13 ( .A1(SubCellInst_SboxInst_13_n8), .A2(
        SubCellInst_SboxInst_13_n7), .ZN(SubCellInst_SboxInst_13_n15) );
  NAND2_X1 SubCellInst_SboxInst_13_U12 ( .A1(SubCellInst_SboxInst_13_n6), .A2(
        SubCellInst_SboxInst_13_n5), .ZN(Feedback[53]) );
  NAND2_X1 SubCellInst_SboxInst_13_U11 ( .A1(ciphertext[8]), .A2(
        SubCellInst_SboxInst_13_n4), .ZN(SubCellInst_SboxInst_13_n5) );
  NAND2_X1 SubCellInst_SboxInst_13_U10 ( .A1(ciphertext[11]), .A2(
        SubCellInst_SboxInst_13_n9), .ZN(SubCellInst_SboxInst_13_n4) );
  NAND2_X1 SubCellInst_SboxInst_13_U9 ( .A1(ciphertext[10]), .A2(
        SubCellInst_SboxInst_13_n8), .ZN(SubCellInst_SboxInst_13_n6) );
  NOR2_X1 SubCellInst_SboxInst_13_U8 ( .A1(SubCellInst_SboxInst_13_n13), .A2(
        SubCellInst_SboxInst_13_n3), .ZN(Feedback[52]) );
  NOR2_X1 SubCellInst_SboxInst_13_U7 ( .A1(ciphertext[9]), .A2(
        SubCellInst_SboxInst_13_n2), .ZN(SubCellInst_SboxInst_13_n3) );
  NOR2_X1 SubCellInst_SboxInst_13_U6 ( .A1(SubCellInst_SboxInst_13_n7), .A2(
        SubCellInst_SboxInst_13_n1), .ZN(SubCellInst_SboxInst_13_n2) );
  NOR2_X1 SubCellInst_SboxInst_13_U5 ( .A1(ciphertext[10]), .A2(ciphertext[11]), .ZN(
        SubCellInst_SboxInst_13_n1) );
  INV_X1 SubCellInst_SboxInst_13_U4 ( .A(ciphertext[8]), .ZN(
        SubCellInst_SboxInst_13_n7) );
  NOR2_X1 SubCellInst_SboxInst_13_U3 ( .A1(SubCellInst_SboxInst_13_n9), .A2(
        SubCellInst_SboxInst_13_n8), .ZN(SubCellInst_SboxInst_13_n13) );
  INV_X1 SubCellInst_SboxInst_13_U2 ( .A(ciphertext[11]), .ZN(
        SubCellInst_SboxInst_13_n8) );
  INV_X1 SubCellInst_SboxInst_13_U1 ( .A(ciphertext[10]), .ZN(
        SubCellInst_SboxInst_13_n9) );
  NAND2_X1 SubCellInst_SboxInst_14_U19 ( .A1(SubCellInst_SboxInst_14_n15), 
        .A2(SubCellInst_SboxInst_14_n14), .ZN(Feedback[59]) );
  OR2_X1 SubCellInst_SboxInst_14_U18 ( .A1(SubCellInst_SboxInst_14_n13), .A2(
        ciphertext[13]), .ZN(SubCellInst_SboxInst_14_n14) );
  NAND2_X1 SubCellInst_SboxInst_14_U17 ( .A1(SubCellInst_SboxInst_14_n15), 
        .A2(SubCellInst_SboxInst_14_n12), .ZN(Feedback[58]) );
  NAND2_X1 SubCellInst_SboxInst_14_U16 ( .A1(SubCellInst_SboxInst_14_n11), 
        .A2(ciphertext[13]), .ZN(SubCellInst_SboxInst_14_n12) );
  NAND2_X1 SubCellInst_SboxInst_14_U15 ( .A1(SubCellInst_SboxInst_14_n10), 
        .A2(SubCellInst_SboxInst_14_n9), .ZN(SubCellInst_SboxInst_14_n11) );
  NAND2_X1 SubCellInst_SboxInst_14_U14 ( .A1(ciphertext[12]), .A2(ciphertext[15]), 
        .ZN(SubCellInst_SboxInst_14_n10) );
  NAND2_X1 SubCellInst_SboxInst_14_U13 ( .A1(SubCellInst_SboxInst_14_n8), .A2(
        SubCellInst_SboxInst_14_n7), .ZN(SubCellInst_SboxInst_14_n15) );
  NAND2_X1 SubCellInst_SboxInst_14_U12 ( .A1(SubCellInst_SboxInst_14_n6), .A2(
        SubCellInst_SboxInst_14_n5), .ZN(Feedback[57]) );
  NAND2_X1 SubCellInst_SboxInst_14_U11 ( .A1(ciphertext[12]), .A2(
        SubCellInst_SboxInst_14_n4), .ZN(SubCellInst_SboxInst_14_n5) );
  NAND2_X1 SubCellInst_SboxInst_14_U10 ( .A1(ciphertext[15]), .A2(
        SubCellInst_SboxInst_14_n9), .ZN(SubCellInst_SboxInst_14_n4) );
  NAND2_X1 SubCellInst_SboxInst_14_U9 ( .A1(ciphertext[14]), .A2(
        SubCellInst_SboxInst_14_n8), .ZN(SubCellInst_SboxInst_14_n6) );
  NOR2_X1 SubCellInst_SboxInst_14_U8 ( .A1(SubCellInst_SboxInst_14_n13), .A2(
        SubCellInst_SboxInst_14_n3), .ZN(Feedback[56]) );
  NOR2_X1 SubCellInst_SboxInst_14_U7 ( .A1(ciphertext[13]), .A2(
        SubCellInst_SboxInst_14_n2), .ZN(SubCellInst_SboxInst_14_n3) );
  NOR2_X1 SubCellInst_SboxInst_14_U6 ( .A1(SubCellInst_SboxInst_14_n7), .A2(
        SubCellInst_SboxInst_14_n1), .ZN(SubCellInst_SboxInst_14_n2) );
  NOR2_X1 SubCellInst_SboxInst_14_U5 ( .A1(ciphertext[14]), .A2(ciphertext[15]), .ZN(
        SubCellInst_SboxInst_14_n1) );
  INV_X1 SubCellInst_SboxInst_14_U4 ( .A(ciphertext[12]), .ZN(
        SubCellInst_SboxInst_14_n7) );
  NOR2_X1 SubCellInst_SboxInst_14_U3 ( .A1(SubCellInst_SboxInst_14_n9), .A2(
        SubCellInst_SboxInst_14_n8), .ZN(SubCellInst_SboxInst_14_n13) );
  INV_X1 SubCellInst_SboxInst_14_U2 ( .A(ciphertext[15]), .ZN(
        SubCellInst_SboxInst_14_n8) );
  INV_X1 SubCellInst_SboxInst_14_U1 ( .A(ciphertext[14]), .ZN(
        SubCellInst_SboxInst_14_n9) );
  NAND2_X1 SubCellInst_SboxInst_15_U19 ( .A1(SubCellInst_SboxInst_15_n15), 
        .A2(SubCellInst_SboxInst_15_n14), .ZN(Feedback[63]) );
  OR2_X1 SubCellInst_SboxInst_15_U18 ( .A1(SubCellInst_SboxInst_15_n13), .A2(
        ciphertext[1]), .ZN(SubCellInst_SboxInst_15_n14) );
  NAND2_X1 SubCellInst_SboxInst_15_U17 ( .A1(SubCellInst_SboxInst_15_n15), 
        .A2(SubCellInst_SboxInst_15_n12), .ZN(Feedback[62]) );
  NAND2_X1 SubCellInst_SboxInst_15_U16 ( .A1(SubCellInst_SboxInst_15_n11), 
        .A2(ciphertext[1]), .ZN(SubCellInst_SboxInst_15_n12) );
  NAND2_X1 SubCellInst_SboxInst_15_U15 ( .A1(SubCellInst_SboxInst_15_n10), 
        .A2(SubCellInst_SboxInst_15_n9), .ZN(SubCellInst_SboxInst_15_n11) );
  NAND2_X1 SubCellInst_SboxInst_15_U14 ( .A1(ciphertext[0]), .A2(ciphertext[3]), .ZN(
        SubCellInst_SboxInst_15_n10) );
  NAND2_X1 SubCellInst_SboxInst_15_U13 ( .A1(SubCellInst_SboxInst_15_n8), .A2(
        SubCellInst_SboxInst_15_n7), .ZN(SubCellInst_SboxInst_15_n15) );
  NAND2_X1 SubCellInst_SboxInst_15_U12 ( .A1(SubCellInst_SboxInst_15_n6), .A2(
        SubCellInst_SboxInst_15_n5), .ZN(Feedback[61]) );
  NAND2_X1 SubCellInst_SboxInst_15_U11 ( .A1(ciphertext[0]), .A2(
        SubCellInst_SboxInst_15_n4), .ZN(SubCellInst_SboxInst_15_n5) );
  NAND2_X1 SubCellInst_SboxInst_15_U10 ( .A1(ciphertext[3]), .A2(
        SubCellInst_SboxInst_15_n9), .ZN(SubCellInst_SboxInst_15_n4) );
  NAND2_X1 SubCellInst_SboxInst_15_U9 ( .A1(ciphertext[2]), .A2(
        SubCellInst_SboxInst_15_n8), .ZN(SubCellInst_SboxInst_15_n6) );
  NOR2_X1 SubCellInst_SboxInst_15_U8 ( .A1(SubCellInst_SboxInst_15_n13), .A2(
        SubCellInst_SboxInst_15_n3), .ZN(Feedback[60]) );
  NOR2_X1 SubCellInst_SboxInst_15_U7 ( .A1(ciphertext[1]), .A2(
        SubCellInst_SboxInst_15_n2), .ZN(SubCellInst_SboxInst_15_n3) );
  NOR2_X1 SubCellInst_SboxInst_15_U6 ( .A1(SubCellInst_SboxInst_15_n7), .A2(
        SubCellInst_SboxInst_15_n1), .ZN(SubCellInst_SboxInst_15_n2) );
  NOR2_X1 SubCellInst_SboxInst_15_U5 ( .A1(ciphertext[2]), .A2(ciphertext[3]), .ZN(
        SubCellInst_SboxInst_15_n1) );
  INV_X1 SubCellInst_SboxInst_15_U4 ( .A(ciphertext[0]), .ZN(
        SubCellInst_SboxInst_15_n7) );
  NOR2_X1 SubCellInst_SboxInst_15_U3 ( .A1(SubCellInst_SboxInst_15_n9), .A2(
        SubCellInst_SboxInst_15_n8), .ZN(SubCellInst_SboxInst_15_n13) );
  INV_X1 SubCellInst_SboxInst_15_U2 ( .A(ciphertext[3]), .ZN(
        SubCellInst_SboxInst_15_n8) );
  INV_X1 SubCellInst_SboxInst_15_U1 ( .A(ciphertext[2]), .ZN(
        SubCellInst_SboxInst_15_n9) );
  INV_X1 KeyMUX_U3 ( .A(selects[0]), .ZN(KeyMUX_n9) );
  INV_X1 KeyMUX_U2 ( .A(KeyMUX_n9), .ZN(KeyMUX_n8) );
  INV_X2 KeyMUX_U1 ( .A(KeyMUX_n9), .ZN(KeyMUX_n7) );
  MUX2_X1 KeyMUX_MUXInst_0_U1 ( .A(key[64]), .B(key[0]), .S(selects[0]), .Z(
        SelectedKey[0]) );
  MUX2_X1 KeyMUX_MUXInst_1_U1 ( .A(key[65]), .B(key[1]), .S(KeyMUX_n8), .Z(
        SelectedKey[1]) );
  MUX2_X1 KeyMUX_MUXInst_2_U1 ( .A(key[66]), .B(key[2]), .S(selects[0]), .Z(
        SelectedKey[2]) );
  MUX2_X1 KeyMUX_MUXInst_3_U1 ( .A(key[67]), .B(key[3]), .S(KeyMUX_n8), .Z(
        SelectedKey[3]) );
  MUX2_X1 KeyMUX_MUXInst_4_U1 ( .A(key[68]), .B(key[4]), .S(KeyMUX_n8), .Z(
        SelectedKey[4]) );
  MUX2_X1 KeyMUX_MUXInst_5_U1 ( .A(key[69]), .B(key[5]), .S(KeyMUX_n8), .Z(
        SelectedKey[5]) );
  MUX2_X1 KeyMUX_MUXInst_6_U1 ( .A(key[70]), .B(key[6]), .S(KeyMUX_n8), .Z(
        SelectedKey[6]) );
  MUX2_X1 KeyMUX_MUXInst_7_U1 ( .A(key[71]), .B(key[7]), .S(KeyMUX_n8), .Z(
        SelectedKey[7]) );
  MUX2_X1 KeyMUX_MUXInst_8_U1 ( .A(key[72]), .B(key[8]), .S(KeyMUX_n8), .Z(
        SelectedKey[8]) );
  MUX2_X1 KeyMUX_MUXInst_9_U1 ( .A(key[73]), .B(key[9]), .S(KeyMUX_n8), .Z(
        SelectedKey[9]) );
  MUX2_X1 KeyMUX_MUXInst_10_U1 ( .A(key[74]), .B(key[10]), .S(KeyMUX_n8), .Z(
        SelectedKey[10]) );
  MUX2_X1 KeyMUX_MUXInst_11_U1 ( .A(key[75]), .B(key[11]), .S(KeyMUX_n8), .Z(
        SelectedKey[11]) );
  MUX2_X1 KeyMUX_MUXInst_12_U1 ( .A(key[76]), .B(key[12]), .S(KeyMUX_n8), .Z(
        SelectedKey[12]) );
  MUX2_X1 KeyMUX_MUXInst_13_U1 ( .A(key[77]), .B(key[13]), .S(KeyMUX_n8), .Z(
        SelectedKey[13]) );
  MUX2_X1 KeyMUX_MUXInst_14_U1 ( .A(key[78]), .B(key[14]), .S(KeyMUX_n8), .Z(
        SelectedKey[14]) );
  MUX2_X1 KeyMUX_MUXInst_15_U1 ( .A(key[79]), .B(key[15]), .S(KeyMUX_n8), .Z(
        SelectedKey[15]) );
  MUX2_X1 KeyMUX_MUXInst_16_U1 ( .A(key[80]), .B(key[16]), .S(KeyMUX_n8), .Z(
        SelectedKey[16]) );
  MUX2_X1 KeyMUX_MUXInst_17_U1 ( .A(key[81]), .B(key[17]), .S(KeyMUX_n8), .Z(
        SelectedKey[17]) );
  MUX2_X1 KeyMUX_MUXInst_18_U1 ( .A(key[82]), .B(key[18]), .S(KeyMUX_n8), .Z(
        SelectedKey[18]) );
  MUX2_X1 KeyMUX_MUXInst_19_U1 ( .A(key[83]), .B(key[19]), .S(KeyMUX_n8), .Z(
        SelectedKey[19]) );
  MUX2_X1 KeyMUX_MUXInst_20_U1 ( .A(key[84]), .B(key[20]), .S(KeyMUX_n8), .Z(
        SelectedKey[20]) );
  MUX2_X1 KeyMUX_MUXInst_21_U1 ( .A(key[85]), .B(key[21]), .S(KeyMUX_n8), .Z(
        SelectedKey[21]) );
  MUX2_X1 KeyMUX_MUXInst_22_U1 ( .A(key[86]), .B(key[22]), .S(selects[0]), .Z(
        SelectedKey[22]) );
  MUX2_X1 KeyMUX_MUXInst_23_U1 ( .A(key[87]), .B(key[23]), .S(selects[0]), .Z(
        SelectedKey[23]) );
  MUX2_X1 KeyMUX_MUXInst_24_U1 ( .A(key[88]), .B(key[24]), .S(selects[0]), .Z(
        SelectedKey[24]) );
  MUX2_X1 KeyMUX_MUXInst_25_U1 ( .A(key[89]), .B(key[25]), .S(selects[0]), .Z(
        SelectedKey[25]) );
  MUX2_X1 KeyMUX_MUXInst_26_U1 ( .A(key[90]), .B(key[26]), .S(selects[0]), .Z(
        SelectedKey[26]) );
  MUX2_X1 KeyMUX_MUXInst_27_U1 ( .A(key[91]), .B(key[27]), .S(selects[0]), .Z(
        SelectedKey[27]) );
  MUX2_X1 KeyMUX_MUXInst_28_U1 ( .A(key[92]), .B(key[28]), .S(KeyMUX_n7), .Z(
        SelectedKey[28]) );
  MUX2_X1 KeyMUX_MUXInst_29_U1 ( .A(key[93]), .B(key[29]), .S(KeyMUX_n7), .Z(
        SelectedKey[29]) );
  MUX2_X1 KeyMUX_MUXInst_30_U1 ( .A(key[94]), .B(key[30]), .S(KeyMUX_n7), .Z(
        SelectedKey[30]) );
  MUX2_X1 KeyMUX_MUXInst_31_U1 ( .A(key[95]), .B(key[31]), .S(KeyMUX_n7), .Z(
        SelectedKey[31]) );
  MUX2_X1 KeyMUX_MUXInst_32_U1 ( .A(key[96]), .B(key[32]), .S(KeyMUX_n7), .Z(
        SelectedKey[32]) );
  MUX2_X1 KeyMUX_MUXInst_33_U1 ( .A(key[97]), .B(key[33]), .S(selects[0]), .Z(
        SelectedKey[33]) );
  MUX2_X1 KeyMUX_MUXInst_34_U1 ( .A(key[98]), .B(key[34]), .S(KeyMUX_n7), .Z(
        SelectedKey[34]) );
  MUX2_X1 KeyMUX_MUXInst_35_U1 ( .A(key[99]), .B(key[35]), .S(KeyMUX_n7), .Z(
        SelectedKey[35]) );
  MUX2_X1 KeyMUX_MUXInst_36_U1 ( .A(key[100]), .B(key[36]), .S(selects[0]), 
        .Z(SelectedKey[36]) );
  MUX2_X1 KeyMUX_MUXInst_37_U1 ( .A(key[101]), .B(key[37]), .S(KeyMUX_n7), .Z(
        SelectedKey[37]) );
  MUX2_X1 KeyMUX_MUXInst_38_U1 ( .A(key[102]), .B(key[38]), .S(KeyMUX_n7), .Z(
        SelectedKey[38]) );
  MUX2_X1 KeyMUX_MUXInst_39_U1 ( .A(key[103]), .B(key[39]), .S(selects[0]), 
        .Z(SelectedKey[39]) );
  MUX2_X1 KeyMUX_MUXInst_40_U1 ( .A(key[104]), .B(key[40]), .S(KeyMUX_n7), .Z(
        SelectedKey[40]) );
  MUX2_X1 KeyMUX_MUXInst_41_U1 ( .A(key[105]), .B(key[41]), .S(KeyMUX_n7), .Z(
        SelectedKey[41]) );
  MUX2_X1 KeyMUX_MUXInst_42_U1 ( .A(key[106]), .B(key[42]), .S(KeyMUX_n7), .Z(
        SelectedKey[42]) );
  MUX2_X1 KeyMUX_MUXInst_43_U1 ( .A(key[107]), .B(key[43]), .S(KeyMUX_n7), .Z(
        SelectedKey[43]) );
  MUX2_X1 KeyMUX_MUXInst_44_U1 ( .A(key[108]), .B(key[44]), .S(KeyMUX_n7), .Z(
        SelectedKey[44]) );
  MUX2_X1 KeyMUX_MUXInst_45_U1 ( .A(key[109]), .B(key[45]), .S(KeyMUX_n7), .Z(
        SelectedKey[45]) );
  MUX2_X1 KeyMUX_MUXInst_46_U1 ( .A(key[110]), .B(key[46]), .S(KeyMUX_n7), .Z(
        SelectedKey[46]) );
  MUX2_X1 KeyMUX_MUXInst_47_U1 ( .A(key[111]), .B(key[47]), .S(KeyMUX_n7), .Z(
        SelectedKey[47]) );
  MUX2_X1 KeyMUX_MUXInst_48_U1 ( .A(key[112]), .B(key[48]), .S(KeyMUX_n7), .Z(
        SelectedKey[48]) );
  MUX2_X1 KeyMUX_MUXInst_49_U1 ( .A(key[113]), .B(key[49]), .S(KeyMUX_n7), .Z(
        SelectedKey[49]) );
  MUX2_X1 KeyMUX_MUXInst_50_U1 ( .A(key[114]), .B(key[50]), .S(KeyMUX_n7), .Z(
        SelectedKey[50]) );
  MUX2_X1 KeyMUX_MUXInst_51_U1 ( .A(key[115]), .B(key[51]), .S(KeyMUX_n7), .Z(
        SelectedKey[51]) );
  MUX2_X1 KeyMUX_MUXInst_52_U1 ( .A(key[116]), .B(key[52]), .S(KeyMUX_n7), .Z(
        SelectedKey[52]) );
  MUX2_X1 KeyMUX_MUXInst_53_U1 ( .A(key[117]), .B(key[53]), .S(selects[0]), 
        .Z(SelectedKey[53]) );
  MUX2_X1 KeyMUX_MUXInst_54_U1 ( .A(key[118]), .B(key[54]), .S(selects[0]), 
        .Z(SelectedKey[54]) );
  MUX2_X1 KeyMUX_MUXInst_55_U1 ( .A(key[119]), .B(key[55]), .S(KeyMUX_n7), .Z(
        SelectedKey[55]) );
  MUX2_X1 KeyMUX_MUXInst_56_U1 ( .A(key[120]), .B(key[56]), .S(selects[0]), 
        .Z(SelectedKey[56]) );
  MUX2_X1 KeyMUX_MUXInst_57_U1 ( .A(key[121]), .B(key[57]), .S(KeyMUX_n7), .Z(
        SelectedKey[57]) );
  MUX2_X1 KeyMUX_MUXInst_58_U1 ( .A(key[122]), .B(key[58]), .S(KeyMUX_n7), .Z(
        SelectedKey[58]) );
  MUX2_X1 KeyMUX_MUXInst_59_U1 ( .A(key[123]), .B(key[59]), .S(selects[0]), 
        .Z(SelectedKey[59]) );
  MUX2_X1 KeyMUX_MUXInst_60_U1 ( .A(key[124]), .B(key[60]), .S(KeyMUX_n7), .Z(
        SelectedKey[60]) );
  MUX2_X1 KeyMUX_MUXInst_61_U1 ( .A(key[125]), .B(key[61]), .S(KeyMUX_n7), .Z(
        SelectedKey[61]) );
  MUX2_X1 KeyMUX_MUXInst_62_U1 ( .A(key[126]), .B(key[62]), .S(selects[0]), 
        .Z(SelectedKey[62]) );
  MUX2_X1 KeyMUX_MUXInst_63_U1 ( .A(key[127]), .B(key[63]), .S(KeyMUX_n7), .Z(
        SelectedKey[63]) );
  MUX2_X1 FSMMUX_MUXInst_0_U1 ( .A(FSMReg[0]), .B(1'b1), .S(rst), .Z(
        RoundConstant_0) );
  MUX2_X1 FSMMUX_MUXInst_1_U1 ( .A(FSMReg[1]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[0]) );
  MUX2_X1 FSMMUX_MUXInst_2_U1 ( .A(FSMReg[2]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[1]) );
  MUX2_X1 FSMMUX_MUXInst_3_U1 ( .A(FSMReg[3]), .B(1'b1), .S(rst), .Z(
        RoundConstant_4_) );
  MUX2_X1 FSMMUX_MUXInst_4_U1 ( .A(FSMReg[4]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[3]) );
  MUX2_X1 FSMMUX_MUXInst_5_U1 ( .A(FSMReg[5]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[4]) );
  MUX2_X1 FSMMUX_MUXInst_6_U1 ( .A(FSMReg[6]), .B(1'b0), .S(rst), .Z(
        FSMUpdate[5]) );
  XOR2_X1 FSMUpdateInst_U2 ( .A(RoundConstant_4_), .B(FSMUpdate[3]), .Z(
        FSMUpdate[6]) );
  XOR2_X1 FSMUpdateInst_U1 ( .A(FSMUpdate[0]), .B(RoundConstant_0), .Z(
        FSMUpdate[2]) );
  INV_X1 FSMRegInst_s_current_state_reg_6__U1 ( .A(FSMReg[6]), .ZN(
        FSMRegInst_s_current_state_reg_6__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_6__FF_FF ( .D(FSMUpdate[6]), .CK(clk), 
        .Q(FSMReg[6]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_5__U1 ( .A(FSMReg[5]), .ZN(
        FSMRegInst_s_current_state_reg_5__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_5__FF_FF ( .D(FSMUpdate[5]), .CK(clk), 
        .Q(FSMReg[5]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_4__U1 ( .A(FSMReg[4]), .ZN(
        FSMRegInst_s_current_state_reg_4__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_4__FF_FF ( .D(FSMUpdate[4]), .CK(clk), 
        .Q(FSMReg[4]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_3__U1 ( .A(FSMReg[3]), .ZN(
        FSMRegInst_s_current_state_reg_3__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_3__FF_FF ( .D(FSMUpdate[3]), .CK(clk), 
        .Q(FSMReg[3]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_2__U1 ( .A(FSMReg[2]), .ZN(
        FSMRegInst_s_current_state_reg_2__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_2__FF_FF ( .D(FSMUpdate[2]), .CK(clk), 
        .Q(FSMReg[2]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_1__U1 ( .A(FSMReg[1]), .ZN(
        FSMRegInst_s_current_state_reg_1__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_1__FF_FF ( .D(FSMUpdate[1]), .CK(clk), 
        .Q(FSMReg[1]), .QN() );
  INV_X1 FSMRegInst_s_current_state_reg_0__U1 ( .A(FSMReg[0]), .ZN(
        FSMRegInst_s_current_state_reg_0__QN) );
  DFF_X1 FSMRegInst_s_current_state_reg_0__FF_FF ( .D(FSMUpdate[0]), .CK(clk), 
        .Q(FSMReg[0]), .QN() );
  AND2_X1 FSMSignalsInst_U6 ( .A1(FSMUpdate[5]), .A2(FSMSignalsInst_n5), .ZN(
        done_internal) );
  NOR2_X1 FSMSignalsInst_U5 ( .A1(FSMSignalsInst_n4), .A2(FSMSignalsInst_n3), 
        .ZN(FSMSignalsInst_n5) );
  NAND2_X1 FSMSignalsInst_U4 ( .A1(FSMSignalsInst_n2), .A2(FSMSignalsInst_n1), 
        .ZN(FSMSignalsInst_n3) );
  NOR2_X1 FSMSignalsInst_U3 ( .A1(FSMUpdate[3]), .A2(FSMUpdate[4]), .ZN(
        FSMSignalsInst_n1) );
  NOR2_X1 FSMSignalsInst_U2 ( .A1(FSMUpdate[0]), .A2(RoundConstant_4_), .ZN(
        FSMSignalsInst_n2) );
  NAND2_X1 FSMSignalsInst_U1 ( .A1(RoundConstant_0), .A2(FSMUpdate[1]), .ZN(
        FSMSignalsInst_n4) );
  MUX2_X1 selectsMUX_MUXInst_0_U1 ( .A(selectsReg[0]), .B(1'b0), .S(rst), .Z(
        selects[0]) );
  MUX2_X1 selectsMUX_MUXInst_1_U1 ( .A(selectsReg[1]), .B(1'b0), .S(rst), .Z(
        selects[1]) );
  XNOR2_X1 selectsUpdateInst_U3 ( .A(selectsUpdateInst_n3), .B(selects[1]), 
        .ZN(selectsNext[1]) );
  XNOR2_X1 selectsUpdateInst_U2 ( .A(selects[0]), .B(1'b0), .ZN(
        selectsUpdateInst_n3) );
  INV_X1 selectsUpdateInst_U1 ( .A(selects[0]), .ZN(selectsNext[0]) );
  INV_X1 selectsRegInst_s_current_state_reg_1__U1 ( .A(selectsReg[1]), .ZN(
        selectsRegInst_s_current_state_reg_1__QN) );
  DFF_X1 selectsRegInst_s_current_state_reg_1__FF_FF ( .D(selectsNext[1]), 
        .CK(clk), .Q(selectsReg[1]), .QN() );
  INV_X1 selectsRegInst_s_current_state_reg_0__U1 ( .A(selectsReg[0]), .ZN(
        selectsRegInst_s_current_state_reg_0__QN) );
  DFF_X1 selectsRegInst_s_current_state_reg_0__FF_FF ( .D(selectsNext[0]), 
        .CK(clk), .Q(selectsReg[0]), .QN() );
  INV_X1 done_reg_U1 ( .A(done), .ZN(done_reg_QN) );
  DFF_X1 done_reg_FF_FF ( .D(done_internal), .CK(clk), .Q(done), .QN() );
endmodule

